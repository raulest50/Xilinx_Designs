

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity stream_source is
    Port (
    clk : in std_logic;
    nrst : in std_logic;
    axis_mtr_tready : in std_logic;
    axis_mtr_tvalid : out std_logic;
    axis_mtr_tdata : out std_logic_vector(12 downto 0)
    );
end stream_source;

architecture Behavioral of stream_source is

type estado is (init, tvalid, tready);
signal n : integer range 0 to 8191 := 0;

type data_8x32 is array (0 to 8191) of std_logic_vector(12 downto 0);

constant my_data : data_8x32  :=
(
     0 => b"0000000000000",  1 => b"0000000000001",  2 => b"0000000000010",  3 => b"0000000000011",
 4 => b"0000000000100",  5 => b"0000000000101",  6 => b"0000000000111",  7 => b"0000000001000",
 8 => b"0000000001001",  9 => b"0000000001010",  10 => b"0000000001011",  11 => b"0000000001100",
 12 => b"0000000001110",  13 => b"0000000001111",  14 => b"0000000010000",  15 => b"0000000010001",
 16 => b"0000000010010",  17 => b"0000000010100",  18 => b"0000000010101",  19 => b"0000000010110",
 20 => b"0000000010111",  21 => b"0000000011000",  22 => b"0000000011001",  23 => b"0000000011011",
 24 => b"0000000011100",  25 => b"0000000011101",  26 => b"0000000011110",  27 => b"0000000011111",
 28 => b"0000000100000",  29 => b"0000000100010",  30 => b"0000000100011",  31 => b"0000000100100",
 32 => b"0000000100101",  33 => b"0000000100110",  34 => b"0000000101000",  35 => b"0000000101001",
 36 => b"0000000101010",  37 => b"0000000101011",  38 => b"0000000101100",  39 => b"0000000101101",
 40 => b"0000000101111",  41 => b"0000000110000",  42 => b"0000000110001",  43 => b"0000000110010",
 44 => b"0000000110011",  45 => b"0000000110100",  46 => b"0000000110110",  47 => b"0000000110111",
 48 => b"0000000111000",  49 => b"0000000111001",  50 => b"0000000111010",  51 => b"0000000111100",
 52 => b"0000000111101",  53 => b"0000000111110",  54 => b"0000000111111",  55 => b"0000001000000",
 56 => b"0000001000001",  57 => b"0000001000011",  58 => b"0000001000100",  59 => b"0000001000101",
 60 => b"0000001000110",  61 => b"0000001000111",  62 => b"0000001001000",  63 => b"0000001001010",
 64 => b"0000001001011",  65 => b"0000001001100",  66 => b"0000001001101",  67 => b"0000001001110",
 68 => b"0000001010000",  69 => b"0000001010001",  70 => b"0000001010010",  71 => b"0000001010011",
 72 => b"0000001010100",  73 => b"0000001010101",  74 => b"0000001010111",  75 => b"0000001011000",
 76 => b"0000001011001",  77 => b"0000001011010",  78 => b"0000001011011",  79 => b"0000001011100",
 80 => b"0000001011110",  81 => b"0000001011111",  82 => b"0000001100000",  83 => b"0000001100001",
 84 => b"0000001100010",  85 => b"0000001100011",  86 => b"0000001100101",  87 => b"0000001100110",
 88 => b"0000001100111",  89 => b"0000001101000",  90 => b"0000001101001",  91 => b"0000001101010",
 92 => b"0000001101100",  93 => b"0000001101101",  94 => b"0000001101110",  95 => b"0000001101111",
 96 => b"0000001110000",  97 => b"0000001110001",  98 => b"0000001110011",  99 => b"0000001110100",
 100 => b"0000001110101",  101 => b"0000001110110",  102 => b"0000001110111",  103 => b"0000001111000",
 104 => b"0000001111010",  105 => b"0000001111011",  106 => b"0000001111100",  107 => b"0000001111101",
 108 => b"0000001111110",  109 => b"0000001111111",  110 => b"0000010000001",  111 => b"0000010000010",
 112 => b"0000010000011",  113 => b"0000010000100",  114 => b"0000010000101",  115 => b"0000010000110",
 116 => b"0000010001000",  117 => b"0000010001001",  118 => b"0000010001010",  119 => b"0000010001011",
 120 => b"0000010001100",  121 => b"0000010001101",  122 => b"0000010001111",  123 => b"0000010010000",
 124 => b"0000010010001",  125 => b"0000010010010",  126 => b"0000010010011",  127 => b"0000010010100",
 128 => b"0000010010110",  129 => b"0000010010111",  130 => b"0000010011000",  131 => b"0000010011001",
 132 => b"0000010011010",  133 => b"0000010011011",  134 => b"0000010011101",  135 => b"0000010011110",
 136 => b"0000010011111",  137 => b"0000010100000",  138 => b"0000010100001",  139 => b"0000010100010",
 140 => b"0000010100100",  141 => b"0000010100101",  142 => b"0000010100110",  143 => b"0000010100111",
 144 => b"0000010101000",  145 => b"0000010101001",  146 => b"0000010101010",  147 => b"0000010101100",
 148 => b"0000010101101",  149 => b"0000010101110",  150 => b"0000010101111",  151 => b"0000010110000",
 152 => b"0000010110001",  153 => b"0000010110011",  154 => b"0000010110100",  155 => b"0000010110101",
 156 => b"0000010110110",  157 => b"0000010110111",  158 => b"0000010111000",  159 => b"0000010111001",
 160 => b"0000010111011",  161 => b"0000010111100",  162 => b"0000010111101",  163 => b"0000010111110",
 164 => b"0000010111111",  165 => b"0000011000000",  166 => b"0000011000010",  167 => b"0000011000011",
 168 => b"0000011000100",  169 => b"0000011000101",  170 => b"0000011000110",  171 => b"0000011000111",
 172 => b"0000011001000",  173 => b"0000011001010",  174 => b"0000011001011",  175 => b"0000011001100",
 176 => b"0000011001101",  177 => b"0000011001110",  178 => b"0000011001111",  179 => b"0000011010000",
 180 => b"0000011010010",  181 => b"0000011010011",  182 => b"0000011010100",  183 => b"0000011010101",
 184 => b"0000011010110",  185 => b"0000011010111",  186 => b"0000011011000",  187 => b"0000011011010",
 188 => b"0000011011011",  189 => b"0000011011100",  190 => b"0000011011101",  191 => b"0000011011110",
 192 => b"0000011011111",  193 => b"0000011100000",  194 => b"0000011100010",  195 => b"0000011100011",
 196 => b"0000011100100",  197 => b"0000011100101",  198 => b"0000011100110",  199 => b"0000011100111",
 200 => b"0000011101000",  201 => b"0000011101010",  202 => b"0000011101011",  203 => b"0000011101100",
 204 => b"0000011101101",  205 => b"0000011101110",  206 => b"0000011101111",  207 => b"0000011110000",
 208 => b"0000011110001",  209 => b"0000011110011",  210 => b"0000011110100",  211 => b"0000011110101",
 212 => b"0000011110110",  213 => b"0000011110111",  214 => b"0000011111000",  215 => b"0000011111001",
 216 => b"0000011111011",  217 => b"0000011111100",  218 => b"0000011111101",  219 => b"0000011111110",
 220 => b"0000011111111",  221 => b"0000100000000",  222 => b"0000100000001",  223 => b"0000100000010",
 224 => b"0000100000100",  225 => b"0000100000101",  226 => b"0000100000110",  227 => b"0000100000111",
 228 => b"0000100001000",  229 => b"0000100001001",  230 => b"0000100001010",  231 => b"0000100001011",
 232 => b"0000100001101",  233 => b"0000100001110",  234 => b"0000100001111",  235 => b"0000100010000",
 236 => b"0000100010001",  237 => b"0000100010010",  238 => b"0000100010011",  239 => b"0000100010100",
 240 => b"0000100010110",  241 => b"0000100010111",  242 => b"0000100011000",  243 => b"0000100011001",
 244 => b"0000100011010",  245 => b"0000100011011",  246 => b"0000100011100",  247 => b"0000100011101",
 248 => b"0000100011110",  249 => b"0000100100000",  250 => b"0000100100001",  251 => b"0000100100010",
 252 => b"0000100100011",  253 => b"0000100100100",  254 => b"0000100100101",  255 => b"0000100100110",
 256 => b"0000100100111",  257 => b"0000100101000",  258 => b"0000100101010",  259 => b"0000100101011",
 260 => b"0000100101100",  261 => b"0000100101101",  262 => b"0000100101110",  263 => b"0000100101111",
 264 => b"0000100110000",  265 => b"0000100110001",  266 => b"0000100110010",  267 => b"0000100110100",
 268 => b"0000100110101",  269 => b"0000100110110",  270 => b"0000100110111",  271 => b"0000100111000",
 272 => b"0000100111001",  273 => b"0000100111010",  274 => b"0000100111011",  275 => b"0000100111100",
 276 => b"0000100111101",  277 => b"0000100111111",  278 => b"0000101000000",  279 => b"0000101000001",
 280 => b"0000101000010",  281 => b"0000101000011",  282 => b"0000101000100",  283 => b"0000101000101",
 284 => b"0000101000110",  285 => b"0000101000111",  286 => b"0000101001000",  287 => b"0000101001010",
 288 => b"0000101001011",  289 => b"0000101001100",  290 => b"0000101001101",  291 => b"0000101001110",
 292 => b"0000101001111",  293 => b"0000101010000",  294 => b"0000101010001",  295 => b"0000101010010",
 296 => b"0000101010011",  297 => b"0000101010100",  298 => b"0000101010110",  299 => b"0000101010111",
 300 => b"0000101011000",  301 => b"0000101011001",  302 => b"0000101011010",  303 => b"0000101011011",
 304 => b"0000101011100",  305 => b"0000101011101",  306 => b"0000101011110",  307 => b"0000101011111",
 308 => b"0000101100000",  309 => b"0000101100001",  310 => b"0000101100011",  311 => b"0000101100100",
 312 => b"0000101100101",  313 => b"0000101100110",  314 => b"0000101100111",  315 => b"0000101101000",
 316 => b"0000101101001",  317 => b"0000101101010",  318 => b"0000101101011",  319 => b"0000101101100",
 320 => b"0000101101101",  321 => b"0000101101110",  322 => b"0000101101111",  323 => b"0000101110001",
 324 => b"0000101110010",  325 => b"0000101110011",  326 => b"0000101110100",  327 => b"0000101110101",
 328 => b"0000101110110",  329 => b"0000101110111",  330 => b"0000101111000",  331 => b"0000101111001",
 332 => b"0000101111010",  333 => b"0000101111011",  334 => b"0000101111100",  335 => b"0000101111101",
 336 => b"0000101111110",  337 => b"0000101111111",  338 => b"0000110000001",  339 => b"0000110000010",
 340 => b"0000110000011",  341 => b"0000110000100",  342 => b"0000110000101",  343 => b"0000110000110",
 344 => b"0000110000111",  345 => b"0000110001000",  346 => b"0000110001001",  347 => b"0000110001010",
 348 => b"0000110001011",  349 => b"0000110001100",  350 => b"0000110001101",  351 => b"0000110001110",
 352 => b"0000110001111",  353 => b"0000110010000",  354 => b"0000110010001",  355 => b"0000110010010",
 356 => b"0000110010100",  357 => b"0000110010101",  358 => b"0000110010110",  359 => b"0000110010111",
 360 => b"0000110011000",  361 => b"0000110011001",  362 => b"0000110011010",  363 => b"0000110011011",
 364 => b"0000110011100",  365 => b"0000110011101",  366 => b"0000110011110",  367 => b"0000110011111",
 368 => b"0000110100000",  369 => b"0000110100001",  370 => b"0000110100010",  371 => b"0000110100011",
 372 => b"0000110100100",  373 => b"0000110100101",  374 => b"0000110100110",  375 => b"0000110100111",
 376 => b"0000110101000",  377 => b"0000110101001",  378 => b"0000110101010",  379 => b"0000110101011",
 380 => b"0000110101101",  381 => b"0000110101110",  382 => b"0000110101111",  383 => b"0000110110000",
 384 => b"0000110110001",  385 => b"0000110110010",  386 => b"0000110110011",  387 => b"0000110110100",
 388 => b"0000110110101",  389 => b"0000110110110",  390 => b"0000110110111",  391 => b"0000110111000",
 392 => b"0000110111001",  393 => b"0000110111010",  394 => b"0000110111011",  395 => b"0000110111100",
 396 => b"0000110111101",  397 => b"0000110111110",  398 => b"0000110111111",  399 => b"0000111000000",
 400 => b"0000111000001",  401 => b"0000111000010",  402 => b"0000111000011",  403 => b"0000111000100",
 404 => b"0000111000101",  405 => b"0000111000110",  406 => b"0000111000111",  407 => b"0000111001000",
 408 => b"0000111001001",  409 => b"0000111001010",  410 => b"0000111001011",  411 => b"0000111001100",
 412 => b"0000111001101",  413 => b"0000111001110",  414 => b"0000111001111",  415 => b"0000111010000",
 416 => b"0000111010001",  417 => b"0000111010010",  418 => b"0000111010011",  419 => b"0000111010100",
 420 => b"0000111010101",  421 => b"0000111010110",  422 => b"0000111010111",  423 => b"0000111011000",
 424 => b"0000111011001",  425 => b"0000111011010",  426 => b"0000111011011",  427 => b"0000111011100",
 428 => b"0000111011101",  429 => b"0000111011110",  430 => b"0000111011111",  431 => b"0000111100000",
 432 => b"0000111100001",  433 => b"0000111100010",  434 => b"0000111100011",  435 => b"0000111100100",
 436 => b"0000111100101",  437 => b"0000111100110",  438 => b"0000111100111",  439 => b"0000111101000",
 440 => b"0000111101001",  441 => b"0000111101010",  442 => b"0000111101011",  443 => b"0000111101100",
 444 => b"0000111101101",  445 => b"0000111101110",  446 => b"0000111101111",  447 => b"0000111110000",
 448 => b"0000111110001",  449 => b"0000111110010",  450 => b"0000111110011",  451 => b"0000111110100",
 452 => b"0000111110101",  453 => b"0000111110110",  454 => b"0000111110111",  455 => b"0000111111000",
 456 => b"0000111111001",  457 => b"0000111111010",  458 => b"0000111111011",  459 => b"0000111111100",
 460 => b"0000111111101",  461 => b"0000111111101",  462 => b"0000111111110",  463 => b"0000111111111",
 464 => b"0001000000000",  465 => b"0001000000001",  466 => b"0001000000010",  467 => b"0001000000011",
 468 => b"0001000000100",  469 => b"0001000000101",  470 => b"0001000000110",  471 => b"0001000000111",
 472 => b"0001000001000",  473 => b"0001000001001",  474 => b"0001000001010",  475 => b"0001000001011",
 476 => b"0001000001100",  477 => b"0001000001101",  478 => b"0001000001110",  479 => b"0001000001111",
 480 => b"0001000010000",  481 => b"0001000010001",  482 => b"0001000010010",  483 => b"0001000010011",
 484 => b"0001000010011",  485 => b"0001000010100",  486 => b"0001000010101",  487 => b"0001000010110",
 488 => b"0001000010111",  489 => b"0001000011000",  490 => b"0001000011001",  491 => b"0001000011010",
 492 => b"0001000011011",  493 => b"0001000011100",  494 => b"0001000011101",  495 => b"0001000011110",
 496 => b"0001000011111",  497 => b"0001000100000",  498 => b"0001000100001",  499 => b"0001000100010",
 500 => b"0001000100010",  501 => b"0001000100011",  502 => b"0001000100100",  503 => b"0001000100101",
 504 => b"0001000100110",  505 => b"0001000100111",  506 => b"0001000101000",  507 => b"0001000101001",
 508 => b"0001000101010",  509 => b"0001000101011",  510 => b"0001000101100",  511 => b"0001000101101",
 512 => b"0001000101110",  513 => b"0001000101110",  514 => b"0001000101111",  515 => b"0001000110000",
 516 => b"0001000110001",  517 => b"0001000110010",  518 => b"0001000110011",  519 => b"0001000110100",
 520 => b"0001000110101",  521 => b"0001000110110",  522 => b"0001000110111",  523 => b"0001000111000",
 524 => b"0001000111000",  525 => b"0001000111001",  526 => b"0001000111010",  527 => b"0001000111011",
 528 => b"0001000111100",  529 => b"0001000111101",  530 => b"0001000111110",  531 => b"0001000111111",
 532 => b"0001001000000",  533 => b"0001001000001",  534 => b"0001001000001",  535 => b"0001001000010",
 536 => b"0001001000011",  537 => b"0001001000100",  538 => b"0001001000101",  539 => b"0001001000110",
 540 => b"0001001000111",  541 => b"0001001001000",  542 => b"0001001001001",  543 => b"0001001001010",
 544 => b"0001001001010",  545 => b"0001001001011",  546 => b"0001001001100",  547 => b"0001001001101",
 548 => b"0001001001110",  549 => b"0001001001111",  550 => b"0001001010000",  551 => b"0001001010001",
 552 => b"0001001010001",  553 => b"0001001010010",  554 => b"0001001010011",  555 => b"0001001010100",
 556 => b"0001001010101",  557 => b"0001001010110",  558 => b"0001001010111",  559 => b"0001001011000",
 560 => b"0001001011000",  561 => b"0001001011001",  562 => b"0001001011010",  563 => b"0001001011011",
 564 => b"0001001011100",  565 => b"0001001011101",  566 => b"0001001011110",  567 => b"0001001011111",
 568 => b"0001001011111",  569 => b"0001001100000",  570 => b"0001001100001",  571 => b"0001001100010",
 572 => b"0001001100011",  573 => b"0001001100100",  574 => b"0001001100101",  575 => b"0001001100101",
 576 => b"0001001100110",  577 => b"0001001100111",  578 => b"0001001101000",  579 => b"0001001101001",
 580 => b"0001001101010",  581 => b"0001001101011",  582 => b"0001001101011",  583 => b"0001001101100",
 584 => b"0001001101101",  585 => b"0001001101110",  586 => b"0001001101111",  587 => b"0001001110000",
 588 => b"0001001110000",  589 => b"0001001110001",  590 => b"0001001110010",  591 => b"0001001110011",
 592 => b"0001001110100",  593 => b"0001001110101",  594 => b"0001001110101",  595 => b"0001001110110",
 596 => b"0001001110111",  597 => b"0001001111000",  598 => b"0001001111001",  599 => b"0001001111010",
 600 => b"0001001111010",  601 => b"0001001111011",  602 => b"0001001111100",  603 => b"0001001111101",
 604 => b"0001001111110",  605 => b"0001001111111",  606 => b"0001001111111",  607 => b"0001010000000",
 608 => b"0001010000001",  609 => b"0001010000010",  610 => b"0001010000011",  611 => b"0001010000011",
 612 => b"0001010000100",  613 => b"0001010000101",  614 => b"0001010000110",  615 => b"0001010000111",
 616 => b"0001010001000",  617 => b"0001010001000",  618 => b"0001010001001",  619 => b"0001010001010",
 620 => b"0001010001011",  621 => b"0001010001100",  622 => b"0001010001100",  623 => b"0001010001101",
 624 => b"0001010001110",  625 => b"0001010001111",  626 => b"0001010010000",  627 => b"0001010010000",
 628 => b"0001010010001",  629 => b"0001010010010",  630 => b"0001010010011",  631 => b"0001010010100",
 632 => b"0001010010100",  633 => b"0001010010101",  634 => b"0001010010110",  635 => b"0001010010111",
 636 => b"0001010010111",  637 => b"0001010011000",  638 => b"0001010011001",  639 => b"0001010011010",
 640 => b"0001010011011",  641 => b"0001010011011",  642 => b"0001010011100",  643 => b"0001010011101",
 644 => b"0001010011110",  645 => b"0001010011111",  646 => b"0001010011111",  647 => b"0001010100000",
 648 => b"0001010100001",  649 => b"0001010100010",  650 => b"0001010100010",  651 => b"0001010100011",
 652 => b"0001010100100",  653 => b"0001010100101",  654 => b"0001010100101",  655 => b"0001010100110",
 656 => b"0001010100111",  657 => b"0001010101000",  658 => b"0001010101001",  659 => b"0001010101001",
 660 => b"0001010101010",  661 => b"0001010101011",  662 => b"0001010101100",  663 => b"0001010101100",
 664 => b"0001010101101",  665 => b"0001010101110",  666 => b"0001010101111",  667 => b"0001010101111",
 668 => b"0001010110000",  669 => b"0001010110001",  670 => b"0001010110010",  671 => b"0001010110010",
 672 => b"0001010110011",  673 => b"0001010110100",  674 => b"0001010110101",  675 => b"0001010110101",
 676 => b"0001010110110",  677 => b"0001010110111",  678 => b"0001010111000",  679 => b"0001010111000",
 680 => b"0001010111001",  681 => b"0001010111010",  682 => b"0001010111010",  683 => b"0001010111011",
 684 => b"0001010111100",  685 => b"0001010111101",  686 => b"0001010111101",  687 => b"0001010111110",
 688 => b"0001010111111",  689 => b"0001011000000",  690 => b"0001011000000",  691 => b"0001011000001",
 692 => b"0001011000010",  693 => b"0001011000010",  694 => b"0001011000011",  695 => b"0001011000100",
 696 => b"0001011000101",  697 => b"0001011000101",  698 => b"0001011000110",  699 => b"0001011000111",
 700 => b"0001011000111",  701 => b"0001011001000",  702 => b"0001011001001",  703 => b"0001011001010",
 704 => b"0001011001010",  705 => b"0001011001011",  706 => b"0001011001100",  707 => b"0001011001100",
 708 => b"0001011001101",  709 => b"0001011001110",  710 => b"0001011001111",  711 => b"0001011001111",
 712 => b"0001011010000",  713 => b"0001011010001",  714 => b"0001011010001",  715 => b"0001011010010",
 716 => b"0001011010011",  717 => b"0001011010011",  718 => b"0001011010100",  719 => b"0001011010101",
 720 => b"0001011010101",  721 => b"0001011010110",  722 => b"0001011010111",  723 => b"0001011011000",
 724 => b"0001011011000",  725 => b"0001011011001",  726 => b"0001011011010",  727 => b"0001011011010",
 728 => b"0001011011011",  729 => b"0001011011100",  730 => b"0001011011100",  731 => b"0001011011101",
 732 => b"0001011011110",  733 => b"0001011011110",  734 => b"0001011011111",  735 => b"0001011100000",
 736 => b"0001011100000",  737 => b"0001011100001",  738 => b"0001011100010",  739 => b"0001011100010",
 740 => b"0001011100011",  741 => b"0001011100100",  742 => b"0001011100100",  743 => b"0001011100101",
 744 => b"0001011100110",  745 => b"0001011100110",  746 => b"0001011100111",  747 => b"0001011101000",
 748 => b"0001011101000",  749 => b"0001011101001",  750 => b"0001011101010",  751 => b"0001011101010",
 752 => b"0001011101011",  753 => b"0001011101011",  754 => b"0001011101100",  755 => b"0001011101101",
 756 => b"0001011101101",  757 => b"0001011101110",  758 => b"0001011101111",  759 => b"0001011101111",
 760 => b"0001011110000",  761 => b"0001011110001",  762 => b"0001011110001",  763 => b"0001011110010",
 764 => b"0001011110011",  765 => b"0001011110011",  766 => b"0001011110100",  767 => b"0001011110100",
 768 => b"0001011110101",  769 => b"0001011110110",  770 => b"0001011110110",  771 => b"0001011110111",
 772 => b"0001011111000",  773 => b"0001011111000",  774 => b"0001011111001",  775 => b"0001011111001",
 776 => b"0001011111010",  777 => b"0001011111011",  778 => b"0001011111011",  779 => b"0001011111100",
 780 => b"0001011111100",  781 => b"0001011111101",  782 => b"0001011111110",  783 => b"0001011111110",
 784 => b"0001011111111",  785 => b"0001100000000",  786 => b"0001100000000",  787 => b"0001100000001",
 788 => b"0001100000001",  789 => b"0001100000010",  790 => b"0001100000011",  791 => b"0001100000011",
 792 => b"0001100000100",  793 => b"0001100000100",  794 => b"0001100000101",  795 => b"0001100000101",
 796 => b"0001100000110",  797 => b"0001100000111",  798 => b"0001100000111",  799 => b"0001100001000",
 800 => b"0001100001000",  801 => b"0001100001001",  802 => b"0001100001010",  803 => b"0001100001010",
 804 => b"0001100001011",  805 => b"0001100001011",  806 => b"0001100001100",  807 => b"0001100001101",
 808 => b"0001100001101",  809 => b"0001100001110",  810 => b"0001100001110",  811 => b"0001100001111",
 812 => b"0001100001111",  813 => b"0001100010000",  814 => b"0001100010001",  815 => b"0001100010001",
 816 => b"0001100010010",  817 => b"0001100010010",  818 => b"0001100010011",  819 => b"0001100010011",
 820 => b"0001100010100",  821 => b"0001100010100",  822 => b"0001100010101",  823 => b"0001100010110",
 824 => b"0001100010110",  825 => b"0001100010111",  826 => b"0001100010111",  827 => b"0001100011000",
 828 => b"0001100011000",  829 => b"0001100011001",  830 => b"0001100011001",  831 => b"0001100011010",
 832 => b"0001100011011",  833 => b"0001100011011",  834 => b"0001100011100",  835 => b"0001100011100",
 836 => b"0001100011101",  837 => b"0001100011101",  838 => b"0001100011110",  839 => b"0001100011110",
 840 => b"0001100011111",  841 => b"0001100011111",  842 => b"0001100100000",  843 => b"0001100100000",
 844 => b"0001100100001",  845 => b"0001100100001",  846 => b"0001100100010",  847 => b"0001100100011",
 848 => b"0001100100011",  849 => b"0001100100100",  850 => b"0001100100100",  851 => b"0001100100101",
 852 => b"0001100100101",  853 => b"0001100100110",  854 => b"0001100100110",  855 => b"0001100100111",
 856 => b"0001100100111",  857 => b"0001100101000",  858 => b"0001100101000",  859 => b"0001100101001",
 860 => b"0001100101001",  861 => b"0001100101010",  862 => b"0001100101010",  863 => b"0001100101011",
 864 => b"0001100101011",  865 => b"0001100101100",  866 => b"0001100101100",  867 => b"0001100101101",
 868 => b"0001100101101",  869 => b"0001100101110",  870 => b"0001100101110",  871 => b"0001100101111",
 872 => b"0001100101111",  873 => b"0001100110000",  874 => b"0001100110000",  875 => b"0001100110001",
 876 => b"0001100110001",  877 => b"0001100110010",  878 => b"0001100110010",  879 => b"0001100110011",
 880 => b"0001100110011",  881 => b"0001100110100",  882 => b"0001100110100",  883 => b"0001100110100",
 884 => b"0001100110101",  885 => b"0001100110101",  886 => b"0001100110110",  887 => b"0001100110110",
 888 => b"0001100110111",  889 => b"0001100110111",  890 => b"0001100111000",  891 => b"0001100111000",
 892 => b"0001100111001",  893 => b"0001100111001",  894 => b"0001100111010",  895 => b"0001100111010",
 896 => b"0001100111011",  897 => b"0001100111011",  898 => b"0001100111011",  899 => b"0001100111100",
 900 => b"0001100111100",  901 => b"0001100111101",  902 => b"0001100111101",  903 => b"0001100111110",
 904 => b"0001100111110",  905 => b"0001100111111",  906 => b"0001100111111",  907 => b"0001100111111",
 908 => b"0001101000000",  909 => b"0001101000000",  910 => b"0001101000001",  911 => b"0001101000001",
 912 => b"0001101000010",  913 => b"0001101000010",  914 => b"0001101000011",  915 => b"0001101000011",
 916 => b"0001101000011",  917 => b"0001101000100",  918 => b"0001101000100",  919 => b"0001101000101",
 920 => b"0001101000101",  921 => b"0001101000110",  922 => b"0001101000110",  923 => b"0001101000110",
 924 => b"0001101000111",  925 => b"0001101000111",  926 => b"0001101001000",  927 => b"0001101001000",
 928 => b"0001101001000",  929 => b"0001101001001",  930 => b"0001101001001",  931 => b"0001101001010",
 932 => b"0001101001010",  933 => b"0001101001010",  934 => b"0001101001011",  935 => b"0001101001011",
 936 => b"0001101001100",  937 => b"0001101001100",  938 => b"0001101001100",  939 => b"0001101001101",
 940 => b"0001101001101",  941 => b"0001101001110",  942 => b"0001101001110",  943 => b"0001101001110",
 944 => b"0001101001111",  945 => b"0001101001111",  946 => b"0001101010000",  947 => b"0001101010000",
 948 => b"0001101010000",  949 => b"0001101010001",  950 => b"0001101010001",  951 => b"0001101010010",
 952 => b"0001101010010",  953 => b"0001101010010",  954 => b"0001101010011",  955 => b"0001101010011",
 956 => b"0001101010011",  957 => b"0001101010100",  958 => b"0001101010100",  959 => b"0001101010101",
 960 => b"0001101010101",  961 => b"0001101010101",  962 => b"0001101010110",  963 => b"0001101010110",
 964 => b"0001101010110",  965 => b"0001101010111",  966 => b"0001101010111",  967 => b"0001101010111",
 968 => b"0001101011000",  969 => b"0001101011000",  970 => b"0001101011001",  971 => b"0001101011001",
 972 => b"0001101011001",  973 => b"0001101011010",  974 => b"0001101011010",  975 => b"0001101011010",
 976 => b"0001101011011",  977 => b"0001101011011",  978 => b"0001101011011",  979 => b"0001101011100",
 980 => b"0001101011100",  981 => b"0001101011100",  982 => b"0001101011101",  983 => b"0001101011101",
 984 => b"0001101011101",  985 => b"0001101011110",  986 => b"0001101011110",  987 => b"0001101011110",
 988 => b"0001101011111",  989 => b"0001101011111",  990 => b"0001101011111",  991 => b"0001101100000",
 992 => b"0001101100000",  993 => b"0001101100000",  994 => b"0001101100001",  995 => b"0001101100001",
 996 => b"0001101100001",  997 => b"0001101100010",  998 => b"0001101100010",  999 => b"0001101100010",
 1000 => b"0001101100011",  1001 => b"0001101100011",  1002 => b"0001101100011",  1003 => b"0001101100011",
 1004 => b"0001101100100",  1005 => b"0001101100100",  1006 => b"0001101100100",  1007 => b"0001101100101",
 1008 => b"0001101100101",  1009 => b"0001101100101",  1010 => b"0001101100110",  1011 => b"0001101100110",
 1012 => b"0001101100110",  1013 => b"0001101100110",  1014 => b"0001101100111",  1015 => b"0001101100111",
 1016 => b"0001101100111",  1017 => b"0001101101000",  1018 => b"0001101101000",  1019 => b"0001101101000",
 1020 => b"0001101101000",  1021 => b"0001101101001",  1022 => b"0001101101001",  1023 => b"0001101101001",
 1024 => b"0001101101010",  1025 => b"0001101101010",  1026 => b"0001101101010",  1027 => b"0001101101010",
 1028 => b"0001101101011",  1029 => b"0001101101011",  1030 => b"0001101101011",  1031 => b"0001101101011",
 1032 => b"0001101101100",  1033 => b"0001101101100",  1034 => b"0001101101100",  1035 => b"0001101101101",
 1036 => b"0001101101101",  1037 => b"0001101101101",  1038 => b"0001101101101",  1039 => b"0001101101110",
 1040 => b"0001101101110",  1041 => b"0001101101110",  1042 => b"0001101101110",  1043 => b"0001101101111",
 1044 => b"0001101101111",  1045 => b"0001101101111",  1046 => b"0001101101111",  1047 => b"0001101110000",
 1048 => b"0001101110000",  1049 => b"0001101110000",  1050 => b"0001101110000",  1051 => b"0001101110001",
 1052 => b"0001101110001",  1053 => b"0001101110001",  1054 => b"0001101110001",  1055 => b"0001101110001",
 1056 => b"0001101110010",  1057 => b"0001101110010",  1058 => b"0001101110010",  1059 => b"0001101110010",
 1060 => b"0001101110011",  1061 => b"0001101110011",  1062 => b"0001101110011",  1063 => b"0001101110011",
 1064 => b"0001101110100",  1065 => b"0001101110100",  1066 => b"0001101110100",  1067 => b"0001101110100",
 1068 => b"0001101110100",  1069 => b"0001101110101",  1070 => b"0001101110101",  1071 => b"0001101110101",
 1072 => b"0001101110101",  1073 => b"0001101110101",  1074 => b"0001101110110",  1075 => b"0001101110110",
 1076 => b"0001101110110",  1077 => b"0001101110110",  1078 => b"0001101110110",  1079 => b"0001101110111",
 1080 => b"0001101110111",  1081 => b"0001101110111",  1082 => b"0001101110111",  1083 => b"0001101110111",
 1084 => b"0001101111000",  1085 => b"0001101111000",  1086 => b"0001101111000",  1087 => b"0001101111000",
 1088 => b"0001101111000",  1089 => b"0001101111001",  1090 => b"0001101111001",  1091 => b"0001101111001",
 1092 => b"0001101111001",  1093 => b"0001101111001",  1094 => b"0001101111010",  1095 => b"0001101111010",
 1096 => b"0001101111010",  1097 => b"0001101111010",  1098 => b"0001101111010",  1099 => b"0001101111010",
 1100 => b"0001101111011",  1101 => b"0001101111011",  1102 => b"0001101111011",  1103 => b"0001101111011",
 1104 => b"0001101111011",  1105 => b"0001101111011",  1106 => b"0001101111100",  1107 => b"0001101111100",
 1108 => b"0001101111100",  1109 => b"0001101111100",  1110 => b"0001101111100",  1111 => b"0001101111100",
 1112 => b"0001101111100",  1113 => b"0001101111101",  1114 => b"0001101111101",  1115 => b"0001101111101",
 1116 => b"0001101111101",  1117 => b"0001101111101",  1118 => b"0001101111101",  1119 => b"0001101111110",
 1120 => b"0001101111110",  1121 => b"0001101111110",  1122 => b"0001101111110",  1123 => b"0001101111110",
 1124 => b"0001101111110",  1125 => b"0001101111110",  1126 => b"0001101111110",  1127 => b"0001101111111",
 1128 => b"0001101111111",  1129 => b"0001101111111",  1130 => b"0001101111111",  1131 => b"0001101111111",
 1132 => b"0001101111111",  1133 => b"0001101111111",  1134 => b"0001110000000",  1135 => b"0001110000000",
 1136 => b"0001110000000",  1137 => b"0001110000000",  1138 => b"0001110000000",  1139 => b"0001110000000",
 1140 => b"0001110000000",  1141 => b"0001110000000",  1142 => b"0001110000000",  1143 => b"0001110000001",
 1144 => b"0001110000001",  1145 => b"0001110000001",  1146 => b"0001110000001",  1147 => b"0001110000001",
 1148 => b"0001110000001",  1149 => b"0001110000001",  1150 => b"0001110000001",  1151 => b"0001110000001",
 1152 => b"0001110000001",  1153 => b"0001110000010",  1154 => b"0001110000010",  1155 => b"0001110000010",
 1156 => b"0001110000010",  1157 => b"0001110000010",  1158 => b"0001110000010",  1159 => b"0001110000010",
 1160 => b"0001110000010",  1161 => b"0001110000010",  1162 => b"0001110000010",  1163 => b"0001110000010",
 1164 => b"0001110000011",  1165 => b"0001110000011",  1166 => b"0001110000011",  1167 => b"0001110000011",
 1168 => b"0001110000011",  1169 => b"0001110000011",  1170 => b"0001110000011",  1171 => b"0001110000011",
 1172 => b"0001110000011",  1173 => b"0001110000011",  1174 => b"0001110000011",  1175 => b"0001110000011",
 1176 => b"0001110000011",  1177 => b"0001110000011",  1178 => b"0001110000011",  1179 => b"0001110000100",
 1180 => b"0001110000100",  1181 => b"0001110000100",  1182 => b"0001110000100",  1183 => b"0001110000100",
 1184 => b"0001110000100",  1185 => b"0001110000100",  1186 => b"0001110000100",  1187 => b"0001110000100",
 1188 => b"0001110000100",  1189 => b"0001110000100",  1190 => b"0001110000100",  1191 => b"0001110000100",
 1192 => b"0001110000100",  1193 => b"0001110000100",  1194 => b"0001110000100",  1195 => b"0001110000100",
 1196 => b"0001110000100",  1197 => b"0001110000100",  1198 => b"0001110000100",  1199 => b"0001110000100",
 1200 => b"0001110000100",  1201 => b"0001110000100",  1202 => b"0001110000100",  1203 => b"0001110000101",
 1204 => b"0001110000101",  1205 => b"0001110000101",  1206 => b"0001110000101",  1207 => b"0001110000101",
 1208 => b"0001110000101",  1209 => b"0001110000101",  1210 => b"0001110000101",  1211 => b"0001110000101",
 1212 => b"0001110000101",  1213 => b"0001110000101",  1214 => b"0001110000101",  1215 => b"0001110000101",
 1216 => b"0001110000101",  1217 => b"0001110000101",  1218 => b"0001110000101",  1219 => b"0001110000101",
 1220 => b"0001110000101",  1221 => b"0001110000101",  1222 => b"0001110000101",  1223 => b"0001110000101",
 1224 => b"0001110000101",  1225 => b"0001110000101",  1226 => b"0001110000101",  1227 => b"0001110000101",
 1228 => b"0001110000101",  1229 => b"0001110000101",  1230 => b"0001110000101",  1231 => b"0001110000101",
 1232 => b"0001110000101",  1233 => b"0001110000101",  1234 => b"0001110000101",  1235 => b"0001110000101",
 1236 => b"0001110000101",  1237 => b"0001110000101",  1238 => b"0001110000100",  1239 => b"0001110000100",
 1240 => b"0001110000100",  1241 => b"0001110000100",  1242 => b"0001110000100",  1243 => b"0001110000100",
 1244 => b"0001110000100",  1245 => b"0001110000100",  1246 => b"0001110000100",  1247 => b"0001110000100",
 1248 => b"0001110000100",  1249 => b"0001110000100",  1250 => b"0001110000100",  1251 => b"0001110000100",
 1252 => b"0001110000100",  1253 => b"0001110000100",  1254 => b"0001110000100",  1255 => b"0001110000100",
 1256 => b"0001110000100",  1257 => b"0001110000100",  1258 => b"0001110000100",  1259 => b"0001110000100",
 1260 => b"0001110000100",  1261 => b"0001110000100",  1262 => b"0001110000011",  1263 => b"0001110000011",
 1264 => b"0001110000011",  1265 => b"0001110000011",  1266 => b"0001110000011",  1267 => b"0001110000011",
 1268 => b"0001110000011",  1269 => b"0001110000011",  1270 => b"0001110000011",  1271 => b"0001110000011",
 1272 => b"0001110000011",  1273 => b"0001110000011",  1274 => b"0001110000011",  1275 => b"0001110000011",
 1276 => b"0001110000011",  1277 => b"0001110000010",  1278 => b"0001110000010",  1279 => b"0001110000010",
 1280 => b"0001110000010",  1281 => b"0001110000010",  1282 => b"0001110000010",  1283 => b"0001110000010",
 1284 => b"0001110000010",  1285 => b"0001110000010",  1286 => b"0001110000010",  1287 => b"0001110000010",
 1288 => b"0001110000010",  1289 => b"0001110000001",  1290 => b"0001110000001",  1291 => b"0001110000001",
 1292 => b"0001110000001",  1293 => b"0001110000001",  1294 => b"0001110000001",  1295 => b"0001110000001",
 1296 => b"0001110000001",  1297 => b"0001110000001",  1298 => b"0001110000001",  1299 => b"0001110000000",
 1300 => b"0001110000000",  1301 => b"0001110000000",  1302 => b"0001110000000",  1303 => b"0001110000000",
 1304 => b"0001110000000",  1305 => b"0001110000000",  1306 => b"0001110000000",  1307 => b"0001110000000",
 1308 => b"0001101111111",  1309 => b"0001101111111",  1310 => b"0001101111111",  1311 => b"0001101111111",
 1312 => b"0001101111111",  1313 => b"0001101111111",  1314 => b"0001101111111",  1315 => b"0001101111111",
 1316 => b"0001101111110",  1317 => b"0001101111110",  1318 => b"0001101111110",  1319 => b"0001101111110",
 1320 => b"0001101111110",  1321 => b"0001101111110",  1322 => b"0001101111110",  1323 => b"0001101111101",
 1324 => b"0001101111101",  1325 => b"0001101111101",  1326 => b"0001101111101",  1327 => b"0001101111101",
 1328 => b"0001101111101",  1329 => b"0001101111101",  1330 => b"0001101111100",  1331 => b"0001101111100",
 1332 => b"0001101111100",  1333 => b"0001101111100",  1334 => b"0001101111100",  1335 => b"0001101111100",
 1336 => b"0001101111011",  1337 => b"0001101111011",  1338 => b"0001101111011",  1339 => b"0001101111011",
 1340 => b"0001101111011",  1341 => b"0001101111011",  1342 => b"0001101111011",  1343 => b"0001101111010",
 1344 => b"0001101111010",  1345 => b"0001101111010",  1346 => b"0001101111010",  1347 => b"0001101111010",
 1348 => b"0001101111001",  1349 => b"0001101111001",  1350 => b"0001101111001",  1351 => b"0001101111001",
 1352 => b"0001101111001",  1353 => b"0001101111001",  1354 => b"0001101111000",  1355 => b"0001101111000",
 1356 => b"0001101111000",  1357 => b"0001101111000",  1358 => b"0001101111000",  1359 => b"0001101110111",
 1360 => b"0001101110111",  1361 => b"0001101110111",  1362 => b"0001101110111",  1363 => b"0001101110111",
 1364 => b"0001101110111",  1365 => b"0001101110110",  1366 => b"0001101110110",  1367 => b"0001101110110",
 1368 => b"0001101110110",  1369 => b"0001101110110",  1370 => b"0001101110101",  1371 => b"0001101110101",
 1372 => b"0001101110101",  1373 => b"0001101110101",  1374 => b"0001101110101",  1375 => b"0001101110100",
 1376 => b"0001101110100",  1377 => b"0001101110100",  1378 => b"0001101110100",  1379 => b"0001101110011",
 1380 => b"0001101110011",  1381 => b"0001101110011",  1382 => b"0001101110011",  1383 => b"0001101110011",
 1384 => b"0001101110010",  1385 => b"0001101110010",  1386 => b"0001101110010",  1387 => b"0001101110010",
 1388 => b"0001101110001",  1389 => b"0001101110001",  1390 => b"0001101110001",  1391 => b"0001101110001",
 1392 => b"0001101110001",  1393 => b"0001101110000",  1394 => b"0001101110000",  1395 => b"0001101110000",
 1396 => b"0001101110000",  1397 => b"0001101101111",  1398 => b"0001101101111",  1399 => b"0001101101111",
 1400 => b"0001101101111",  1401 => b"0001101101110",  1402 => b"0001101101110",  1403 => b"0001101101110",
 1404 => b"0001101101110",  1405 => b"0001101101101",  1406 => b"0001101101101",  1407 => b"0001101101101",
 1408 => b"0001101101101",  1409 => b"0001101101100",  1410 => b"0001101101100",  1411 => b"0001101101100",
 1412 => b"0001101101100",  1413 => b"0001101101011",  1414 => b"0001101101011",  1415 => b"0001101101011",
 1416 => b"0001101101011",  1417 => b"0001101101010",  1418 => b"0001101101010",  1419 => b"0001101101010",
 1420 => b"0001101101010",  1421 => b"0001101101001",  1422 => b"0001101101001",  1423 => b"0001101101001",
 1424 => b"0001101101001",  1425 => b"0001101101000",  1426 => b"0001101101000",  1427 => b"0001101101000",
 1428 => b"0001101100111",  1429 => b"0001101100111",  1430 => b"0001101100111",  1431 => b"0001101100111",
 1432 => b"0001101100110",  1433 => b"0001101100110",  1434 => b"0001101100110",  1435 => b"0001101100101",
 1436 => b"0001101100101",  1437 => b"0001101100101",  1438 => b"0001101100101",  1439 => b"0001101100100",
 1440 => b"0001101100100",  1441 => b"0001101100100",  1442 => b"0001101100011",  1443 => b"0001101100011",
 1444 => b"0001101100011",  1445 => b"0001101100011",  1446 => b"0001101100010",  1447 => b"0001101100010",
 1448 => b"0001101100010",  1449 => b"0001101100001",  1450 => b"0001101100001",  1451 => b"0001101100001",
 1452 => b"0001101100000",  1453 => b"0001101100000",  1454 => b"0001101100000",  1455 => b"0001101100000",
 1456 => b"0001101011111",  1457 => b"0001101011111",  1458 => b"0001101011111",  1459 => b"0001101011110",
 1460 => b"0001101011110",  1461 => b"0001101011110",  1462 => b"0001101011101",  1463 => b"0001101011101",
 1464 => b"0001101011101",  1465 => b"0001101011100",  1466 => b"0001101011100",  1467 => b"0001101011100",
 1468 => b"0001101011011",  1469 => b"0001101011011",  1470 => b"0001101011011",  1471 => b"0001101011010",
 1472 => b"0001101011010",  1473 => b"0001101011010",  1474 => b"0001101011001",  1475 => b"0001101011001",
 1476 => b"0001101011001",  1477 => b"0001101011000",  1478 => b"0001101011000",  1479 => b"0001101011000",
 1480 => b"0001101010111",  1481 => b"0001101010111",  1482 => b"0001101010111",  1483 => b"0001101010110",
 1484 => b"0001101010110",  1485 => b"0001101010110",  1486 => b"0001101010101",  1487 => b"0001101010101",
 1488 => b"0001101010101",  1489 => b"0001101010100",  1490 => b"0001101010100",  1491 => b"0001101010100",
 1492 => b"0001101010011",  1493 => b"0001101010011",  1494 => b"0001101010011",  1495 => b"0001101010010",
 1496 => b"0001101010010",  1497 => b"0001101010001",  1498 => b"0001101010001",  1499 => b"0001101010001",
 1500 => b"0001101010000",  1501 => b"0001101010000",  1502 => b"0001101010000",  1503 => b"0001101001111",
 1504 => b"0001101001111",  1505 => b"0001101001111",  1506 => b"0001101001110",  1507 => b"0001101001110",
 1508 => b"0001101001101",  1509 => b"0001101001101",  1510 => b"0001101001101",  1511 => b"0001101001100",
 1512 => b"0001101001100",  1513 => b"0001101001100",  1514 => b"0001101001011",  1515 => b"0001101001011",
 1516 => b"0001101001010",  1517 => b"0001101001010",  1518 => b"0001101001010",  1519 => b"0001101001001",
 1520 => b"0001101001001",  1521 => b"0001101001000",  1522 => b"0001101001000",  1523 => b"0001101001000",
 1524 => b"0001101000111",  1525 => b"0001101000111",  1526 => b"0001101000110",  1527 => b"0001101000110",
 1528 => b"0001101000110",  1529 => b"0001101000101",  1530 => b"0001101000101",  1531 => b"0001101000101",
 1532 => b"0001101000100",  1533 => b"0001101000100",  1534 => b"0001101000011",  1535 => b"0001101000011",
 1536 => b"0001101000010",  1537 => b"0001101000010",  1538 => b"0001101000010",  1539 => b"0001101000001",
 1540 => b"0001101000001",  1541 => b"0001101000000",  1542 => b"0001101000000",  1543 => b"0001101000000",
 1544 => b"0001100111111",  1545 => b"0001100111111",  1546 => b"0001100111110",  1547 => b"0001100111110",
 1548 => b"0001100111110",  1549 => b"0001100111101",  1550 => b"0001100111101",  1551 => b"0001100111100",
 1552 => b"0001100111100",  1553 => b"0001100111011",  1554 => b"0001100111011",  1555 => b"0001100111011",
 1556 => b"0001100111010",  1557 => b"0001100111010",  1558 => b"0001100111001",  1559 => b"0001100111001",
 1560 => b"0001100111000",  1561 => b"0001100111000",  1562 => b"0001100111000",  1563 => b"0001100110111",
 1564 => b"0001100110111",  1565 => b"0001100110110",  1566 => b"0001100110110",  1567 => b"0001100110101",
 1568 => b"0001100110101",  1569 => b"0001100110101",  1570 => b"0001100110100",  1571 => b"0001100110100",
 1572 => b"0001100110011",  1573 => b"0001100110011",  1574 => b"0001100110010",  1575 => b"0001100110010",
 1576 => b"0001100110001",  1577 => b"0001100110001",  1578 => b"0001100110000",  1579 => b"0001100110000",
 1580 => b"0001100110000",  1581 => b"0001100101111",  1582 => b"0001100101111",  1583 => b"0001100101110",
 1584 => b"0001100101110",  1585 => b"0001100101101",  1586 => b"0001100101101",  1587 => b"0001100101100",
 1588 => b"0001100101100",  1589 => b"0001100101011",  1590 => b"0001100101011",  1591 => b"0001100101011",
 1592 => b"0001100101010",  1593 => b"0001100101010",  1594 => b"0001100101001",  1595 => b"0001100101001",
 1596 => b"0001100101000",  1597 => b"0001100101000",  1598 => b"0001100100111",  1599 => b"0001100100111",
 1600 => b"0001100100110",  1601 => b"0001100100110",  1602 => b"0001100100101",  1603 => b"0001100100101",
 1604 => b"0001100100100",  1605 => b"0001100100100",  1606 => b"0001100100011",  1607 => b"0001100100011",
 1608 => b"0001100100010",  1609 => b"0001100100010",  1610 => b"0001100100001",  1611 => b"0001100100001",
 1612 => b"0001100100001",  1613 => b"0001100100000",  1614 => b"0001100100000",  1615 => b"0001100011111",
 1616 => b"0001100011111",  1617 => b"0001100011110",  1618 => b"0001100011110",  1619 => b"0001100011101",
 1620 => b"0001100011101",  1621 => b"0001100011100",  1622 => b"0001100011100",  1623 => b"0001100011011",
 1624 => b"0001100011011",  1625 => b"0001100011010",  1626 => b"0001100011010",  1627 => b"0001100011001",
 1628 => b"0001100011001",  1629 => b"0001100011000",  1630 => b"0001100011000",  1631 => b"0001100010111",
 1632 => b"0001100010111",  1633 => b"0001100010110",  1634 => b"0001100010110",  1635 => b"0001100010101",
 1636 => b"0001100010101",  1637 => b"0001100010100",  1638 => b"0001100010011",  1639 => b"0001100010011",
 1640 => b"0001100010010",  1641 => b"0001100010010",  1642 => b"0001100010001",  1643 => b"0001100010001",
 1644 => b"0001100010000",  1645 => b"0001100010000",  1646 => b"0001100001111",  1647 => b"0001100001111",
 1648 => b"0001100001110",  1649 => b"0001100001110",  1650 => b"0001100001101",  1651 => b"0001100001101",
 1652 => b"0001100001100",  1653 => b"0001100001100",  1654 => b"0001100001011",  1655 => b"0001100001011",
 1656 => b"0001100001010",  1657 => b"0001100001010",  1658 => b"0001100001001",  1659 => b"0001100001000",
 1660 => b"0001100001000",  1661 => b"0001100000111",  1662 => b"0001100000111",  1663 => b"0001100000110",
 1664 => b"0001100000110",  1665 => b"0001100000101",  1666 => b"0001100000101",  1667 => b"0001100000100",
 1668 => b"0001100000100",  1669 => b"0001100000011",  1670 => b"0001100000011",  1671 => b"0001100000010",
 1672 => b"0001100000001",  1673 => b"0001100000001",  1674 => b"0001100000000",  1675 => b"0001100000000",
 1676 => b"0001011111111",  1677 => b"0001011111111",  1678 => b"0001011111110",  1679 => b"0001011111110",
 1680 => b"0001011111101",  1681 => b"0001011111100",  1682 => b"0001011111100",  1683 => b"0001011111011",
 1684 => b"0001011111011",  1685 => b"0001011111010",  1686 => b"0001011111010",  1687 => b"0001011111001",
 1688 => b"0001011111001",  1689 => b"0001011111000",  1690 => b"0001011110111",  1691 => b"0001011110111",
 1692 => b"0001011110110",  1693 => b"0001011110110",  1694 => b"0001011110101",  1695 => b"0001011110101",
 1696 => b"0001011110100",  1697 => b"0001011110011",  1698 => b"0001011110011",  1699 => b"0001011110010",
 1700 => b"0001011110010",  1701 => b"0001011110001",  1702 => b"0001011110001",  1703 => b"0001011110000",
 1704 => b"0001011101111",  1705 => b"0001011101111",  1706 => b"0001011101110",  1707 => b"0001011101110",
 1708 => b"0001011101101",  1709 => b"0001011101101",  1710 => b"0001011101100",  1711 => b"0001011101011",
 1712 => b"0001011101011",  1713 => b"0001011101010",  1714 => b"0001011101010",  1715 => b"0001011101001",
 1716 => b"0001011101000",  1717 => b"0001011101000",  1718 => b"0001011100111",  1719 => b"0001011100111",
 1720 => b"0001011100110",  1721 => b"0001011100110",  1722 => b"0001011100101",  1723 => b"0001011100100",
 1724 => b"0001011100100",  1725 => b"0001011100011",  1726 => b"0001011100011",  1727 => b"0001011100010",
 1728 => b"0001011100001",  1729 => b"0001011100001",  1730 => b"0001011100000",  1731 => b"0001011100000",
 1732 => b"0001011011111",  1733 => b"0001011011110",  1734 => b"0001011011110",  1735 => b"0001011011101",
 1736 => b"0001011011101",  1737 => b"0001011011100",  1738 => b"0001011011011",  1739 => b"0001011011011",
 1740 => b"0001011011010",  1741 => b"0001011011010",  1742 => b"0001011011001",  1743 => b"0001011011000",
 1744 => b"0001011011000",  1745 => b"0001011010111",  1746 => b"0001011010110",  1747 => b"0001011010110",
 1748 => b"0001011010101",  1749 => b"0001011010101",  1750 => b"0001011010100",  1751 => b"0001011010011",
 1752 => b"0001011010011",  1753 => b"0001011010010",  1754 => b"0001011010010",  1755 => b"0001011010001",
 1756 => b"0001011010000",  1757 => b"0001011010000",  1758 => b"0001011001111",  1759 => b"0001011001110",
 1760 => b"0001011001110",  1761 => b"0001011001101",  1762 => b"0001011001101",  1763 => b"0001011001100",
 1764 => b"0001011001011",  1765 => b"0001011001011",  1766 => b"0001011001010",  1767 => b"0001011001001",
 1768 => b"0001011001001",  1769 => b"0001011001000",  1770 => b"0001011001000",  1771 => b"0001011000111",
 1772 => b"0001011000110",  1773 => b"0001011000110",  1774 => b"0001011000101",  1775 => b"0001011000100",
 1776 => b"0001011000100",  1777 => b"0001011000011",  1778 => b"0001011000010",  1779 => b"0001011000010",
 1780 => b"0001011000001",  1781 => b"0001011000001",  1782 => b"0001011000000",  1783 => b"0001010111111",
 1784 => b"0001010111111",  1785 => b"0001010111110",  1786 => b"0001010111101",  1787 => b"0001010111101",
 1788 => b"0001010111100",  1789 => b"0001010111011",  1790 => b"0001010111011",  1791 => b"0001010111010",
 1792 => b"0001010111001",  1793 => b"0001010111001",  1794 => b"0001010111000",  1795 => b"0001010111000",
 1796 => b"0001010110111",  1797 => b"0001010110110",  1798 => b"0001010110110",  1799 => b"0001010110101",
 1800 => b"0001010110100",  1801 => b"0001010110100",  1802 => b"0001010110011",  1803 => b"0001010110010",
 1804 => b"0001010110010",  1805 => b"0001010110001",  1806 => b"0001010110000",  1807 => b"0001010110000",
 1808 => b"0001010101111",  1809 => b"0001010101110",  1810 => b"0001010101110",  1811 => b"0001010101101",
 1812 => b"0001010101100",  1813 => b"0001010101100",  1814 => b"0001010101011",  1815 => b"0001010101010",
 1816 => b"0001010101010",  1817 => b"0001010101001",  1818 => b"0001010101000",  1819 => b"0001010101000",
 1820 => b"0001010100111",  1821 => b"0001010100110",  1822 => b"0001010100110",  1823 => b"0001010100101",
 1824 => b"0001010100100",  1825 => b"0001010100100",  1826 => b"0001010100011",  1827 => b"0001010100010",
 1828 => b"0001010100010",  1829 => b"0001010100001",  1830 => b"0001010100000",  1831 => b"0001010100000",
 1832 => b"0001010011111",  1833 => b"0001010011110",  1834 => b"0001010011110",  1835 => b"0001010011101",
 1836 => b"0001010011100",  1837 => b"0001010011011",  1838 => b"0001010011011",  1839 => b"0001010011010",
 1840 => b"0001010011001",  1841 => b"0001010011001",  1842 => b"0001010011000",  1843 => b"0001010010111",
 1844 => b"0001010010111",  1845 => b"0001010010110",  1846 => b"0001010010101",  1847 => b"0001010010101",
 1848 => b"0001010010100",  1849 => b"0001010010011",  1850 => b"0001010010011",  1851 => b"0001010010010",
 1852 => b"0001010010001",  1853 => b"0001010010001",  1854 => b"0001010010000",  1855 => b"0001010001111",
 1856 => b"0001010001110",  1857 => b"0001010001110",  1858 => b"0001010001101",  1859 => b"0001010001100",
 1860 => b"0001010001100",  1861 => b"0001010001011",  1862 => b"0001010001010",  1863 => b"0001010001010",
 1864 => b"0001010001001",  1865 => b"0001010001000",  1866 => b"0001010000111",  1867 => b"0001010000111",
 1868 => b"0001010000110",  1869 => b"0001010000101",  1870 => b"0001010000101",  1871 => b"0001010000100",
 1872 => b"0001010000011",  1873 => b"0001010000011",  1874 => b"0001010000010",  1875 => b"0001010000001",
 1876 => b"0001010000000",  1877 => b"0001010000000",  1878 => b"0001001111111",  1879 => b"0001001111110",
 1880 => b"0001001111110",  1881 => b"0001001111101",  1882 => b"0001001111100",  1883 => b"0001001111011",
 1884 => b"0001001111011",  1885 => b"0001001111010",  1886 => b"0001001111001",  1887 => b"0001001111001",
 1888 => b"0001001111000",  1889 => b"0001001110111",  1890 => b"0001001110110",  1891 => b"0001001110110",
 1892 => b"0001001110101",  1893 => b"0001001110100",  1894 => b"0001001110100",  1895 => b"0001001110011",
 1896 => b"0001001110010",  1897 => b"0001001110001",  1898 => b"0001001110001",  1899 => b"0001001110000",
 1900 => b"0001001101111",  1901 => b"0001001101111",  1902 => b"0001001101110",  1903 => b"0001001101101",
 1904 => b"0001001101100",  1905 => b"0001001101100",  1906 => b"0001001101011",  1907 => b"0001001101010",
 1908 => b"0001001101001",  1909 => b"0001001101001",  1910 => b"0001001101000",  1911 => b"0001001100111",
 1912 => b"0001001100111",  1913 => b"0001001100110",  1914 => b"0001001100101",  1915 => b"0001001100100",
 1916 => b"0001001100100",  1917 => b"0001001100011",  1918 => b"0001001100010",  1919 => b"0001001100001",
 1920 => b"0001001100001",  1921 => b"0001001100000",  1922 => b"0001001011111",  1923 => b"0001001011111",
 1924 => b"0001001011110",  1925 => b"0001001011101",  1926 => b"0001001011100",  1927 => b"0001001011100",
 1928 => b"0001001011011",  1929 => b"0001001011010",  1930 => b"0001001011001",  1931 => b"0001001011001",
 1932 => b"0001001011000",  1933 => b"0001001010111",  1934 => b"0001001010110",  1935 => b"0001001010110",
 1936 => b"0001001010101",  1937 => b"0001001010100",  1938 => b"0001001010011",  1939 => b"0001001010011",
 1940 => b"0001001010010",  1941 => b"0001001010001",  1942 => b"0001001010001",  1943 => b"0001001010000",
 1944 => b"0001001001111",  1945 => b"0001001001110",  1946 => b"0001001001110",  1947 => b"0001001001101",
 1948 => b"0001001001100",  1949 => b"0001001001011",  1950 => b"0001001001011",  1951 => b"0001001001010",
 1952 => b"0001001001001",  1953 => b"0001001001000",  1954 => b"0001001001000",  1955 => b"0001001000111",
 1956 => b"0001001000110",  1957 => b"0001001000101",  1958 => b"0001001000101",  1959 => b"0001001000100",
 1960 => b"0001001000011",  1961 => b"0001001000010",  1962 => b"0001001000010",  1963 => b"0001001000001",
 1964 => b"0001001000000",  1965 => b"0001000111111",  1966 => b"0001000111111",  1967 => b"0001000111110",
 1968 => b"0001000111101",  1969 => b"0001000111100",  1970 => b"0001000111100",  1971 => b"0001000111011",
 1972 => b"0001000111010",  1973 => b"0001000111001",  1974 => b"0001000111000",  1975 => b"0001000111000",
 1976 => b"0001000110111",  1977 => b"0001000110110",  1978 => b"0001000110101",  1979 => b"0001000110101",
 1980 => b"0001000110100",  1981 => b"0001000110011",  1982 => b"0001000110010",  1983 => b"0001000110010",
 1984 => b"0001000110001",  1985 => b"0001000110000",  1986 => b"0001000101111",  1987 => b"0001000101111",
 1988 => b"0001000101110",  1989 => b"0001000101101",  1990 => b"0001000101100",  1991 => b"0001000101100",
 1992 => b"0001000101011",  1993 => b"0001000101010",  1994 => b"0001000101001",  1995 => b"0001000101000",
 1996 => b"0001000101000",  1997 => b"0001000100111",  1998 => b"0001000100110",  1999 => b"0001000100101",
 2000 => b"0001000100101",  2001 => b"0001000100100",  2002 => b"0001000100011",  2003 => b"0001000100010",
 2004 => b"0001000100010",  2005 => b"0001000100001",  2006 => b"0001000100000",  2007 => b"0001000011111",
 2008 => b"0001000011110",  2009 => b"0001000011110",  2010 => b"0001000011101",  2011 => b"0001000011100",
 2012 => b"0001000011011",  2013 => b"0001000011011",  2014 => b"0001000011010",  2015 => b"0001000011001",
 2016 => b"0001000011000",  2017 => b"0001000011000",  2018 => b"0001000010111",  2019 => b"0001000010110",
 2020 => b"0001000010101",  2021 => b"0001000010100",  2022 => b"0001000010100",  2023 => b"0001000010011",
 2024 => b"0001000010010",  2025 => b"0001000010001",  2026 => b"0001000010001",  2027 => b"0001000010000",
 2028 => b"0001000001111",  2029 => b"0001000001110",  2030 => b"0001000001101",  2031 => b"0001000001101",
 2032 => b"0001000001100",  2033 => b"0001000001011",  2034 => b"0001000001010",  2035 => b"0001000001001",
 2036 => b"0001000001001",  2037 => b"0001000001000",  2038 => b"0001000000111",  2039 => b"0001000000110",
 2040 => b"0001000000110",  2041 => b"0001000000101",  2042 => b"0001000000100",  2043 => b"0001000000011",
 2044 => b"0001000000010",  2045 => b"0001000000010",  2046 => b"0001000000001",  2047 => b"0001000000000",
 2048 => b"0000111111111",  2049 => b"0000111111111",  2050 => b"0000111111110",  2051 => b"0000111111101",
 2052 => b"0000111111100",  2053 => b"0000111111011",  2054 => b"0000111111011",  2055 => b"0000111111010",
 2056 => b"0000111111001",  2057 => b"0000111111000",  2058 => b"0000111110111",  2059 => b"0000111110111",
 2060 => b"0000111110110",  2061 => b"0000111110101",  2062 => b"0000111110100",  2063 => b"0000111110011",
 2064 => b"0000111110011",  2065 => b"0000111110010",  2066 => b"0000111110001",  2067 => b"0000111110000",
 2068 => b"0000111110000",  2069 => b"0000111101111",  2070 => b"0000111101110",  2071 => b"0000111101101",
 2072 => b"0000111101100",  2073 => b"0000111101100",  2074 => b"0000111101011",  2075 => b"0000111101010",
 2076 => b"0000111101001",  2077 => b"0000111101000",  2078 => b"0000111101000",  2079 => b"0000111100111",
 2080 => b"0000111100110",  2081 => b"0000111100101",  2082 => b"0000111100100",  2083 => b"0000111100100",
 2084 => b"0000111100011",  2085 => b"0000111100010",  2086 => b"0000111100001",  2087 => b"0000111100000",
 2088 => b"0000111100000",  2089 => b"0000111011111",  2090 => b"0000111011110",  2091 => b"0000111011101",
 2092 => b"0000111011100",  2093 => b"0000111011100",  2094 => b"0000111011011",  2095 => b"0000111011010",
 2096 => b"0000111011001",  2097 => b"0000111011000",  2098 => b"0000111011000",  2099 => b"0000111010111",
 2100 => b"0000111010110",  2101 => b"0000111010101",  2102 => b"0000111010100",  2103 => b"0000111010100",
 2104 => b"0000111010011",  2105 => b"0000111010010",  2106 => b"0000111010001",  2107 => b"0000111010000",
 2108 => b"0000111010000",  2109 => b"0000111001111",  2110 => b"0000111001110",  2111 => b"0000111001101",
 2112 => b"0000111001100",  2113 => b"0000111001100",  2114 => b"0000111001011",  2115 => b"0000111001010",
 2116 => b"0000111001001",  2117 => b"0000111001000",  2118 => b"0000111001000",  2119 => b"0000111000111",
 2120 => b"0000111000110",  2121 => b"0000111000101",  2122 => b"0000111000100",  2123 => b"0000111000100",
 2124 => b"0000111000011",  2125 => b"0000111000010",  2126 => b"0000111000001",  2127 => b"0000111000000",
 2128 => b"0000111000000",  2129 => b"0000110111111",  2130 => b"0000110111110",  2131 => b"0000110111101",
 2132 => b"0000110111100",  2133 => b"0000110111100",  2134 => b"0000110111011",  2135 => b"0000110111010",
 2136 => b"0000110111001",  2137 => b"0000110111000",  2138 => b"0000110111000",  2139 => b"0000110110111",
 2140 => b"0000110110110",  2141 => b"0000110110101",  2142 => b"0000110110100",  2143 => b"0000110110100",
 2144 => b"0000110110011",  2145 => b"0000110110010",  2146 => b"0000110110001",  2147 => b"0000110110000",
 2148 => b"0000110110000",  2149 => b"0000110101111",  2150 => b"0000110101110",  2151 => b"0000110101101",
 2152 => b"0000110101100",  2153 => b"0000110101100",  2154 => b"0000110101011",  2155 => b"0000110101010",
 2156 => b"0000110101001",  2157 => b"0000110101000",  2158 => b"0000110100111",  2159 => b"0000110100111",
 2160 => b"0000110100110",  2161 => b"0000110100101",  2162 => b"0000110100100",  2163 => b"0000110100011",
 2164 => b"0000110100011",  2165 => b"0000110100010",  2166 => b"0000110100001",  2167 => b"0000110100000",
 2168 => b"0000110011111",  2169 => b"0000110011111",  2170 => b"0000110011110",  2171 => b"0000110011101",
 2172 => b"0000110011100",  2173 => b"0000110011011",  2174 => b"0000110011011",  2175 => b"0000110011010",
 2176 => b"0000110011001",  2177 => b"0000110011000",  2178 => b"0000110010111",  2179 => b"0000110010111",
 2180 => b"0000110010110",  2181 => b"0000110010101",  2182 => b"0000110010100",  2183 => b"0000110010011",
 2184 => b"0000110010010",  2185 => b"0000110010010",  2186 => b"0000110010001",  2187 => b"0000110010000",
 2188 => b"0000110001111",  2189 => b"0000110001110",  2190 => b"0000110001110",  2191 => b"0000110001101",
 2192 => b"0000110001100",  2193 => b"0000110001011",  2194 => b"0000110001010",  2195 => b"0000110001010",
 2196 => b"0000110001001",  2197 => b"0000110001000",  2198 => b"0000110000111",  2199 => b"0000110000110",
 2200 => b"0000110000110",  2201 => b"0000110000101",  2202 => b"0000110000100",  2203 => b"0000110000011",
 2204 => b"0000110000010",  2205 => b"0000110000001",  2206 => b"0000110000001",  2207 => b"0000110000000",
 2208 => b"0000101111111",  2209 => b"0000101111110",  2210 => b"0000101111101",  2211 => b"0000101111101",
 2212 => b"0000101111100",  2213 => b"0000101111011",  2214 => b"0000101111010",  2215 => b"0000101111001",
 2216 => b"0000101111001",  2217 => b"0000101111000",  2218 => b"0000101110111",  2219 => b"0000101110110",
 2220 => b"0000101110101",  2221 => b"0000101110100",  2222 => b"0000101110100",  2223 => b"0000101110011",
 2224 => b"0000101110010",  2225 => b"0000101110001",  2226 => b"0000101110000",  2227 => b"0000101110000",
 2228 => b"0000101101111",  2229 => b"0000101101110",  2230 => b"0000101101101",  2231 => b"0000101101100",
 2232 => b"0000101101100",  2233 => b"0000101101011",  2234 => b"0000101101010",  2235 => b"0000101101001",
 2236 => b"0000101101000",  2237 => b"0000101101000",  2238 => b"0000101100111",  2239 => b"0000101100110",
 2240 => b"0000101100101",  2241 => b"0000101100100",  2242 => b"0000101100011",  2243 => b"0000101100011",
 2244 => b"0000101100010",  2245 => b"0000101100001",  2246 => b"0000101100000",  2247 => b"0000101011111",
 2248 => b"0000101011111",  2249 => b"0000101011110",  2250 => b"0000101011101",  2251 => b"0000101011100",
 2252 => b"0000101011011",  2253 => b"0000101011011",  2254 => b"0000101011010",  2255 => b"0000101011001",
 2256 => b"0000101011000",  2257 => b"0000101010111",  2258 => b"0000101010111",  2259 => b"0000101010110",
 2260 => b"0000101010101",  2261 => b"0000101010100",  2262 => b"0000101010011",  2263 => b"0000101010011",
 2264 => b"0000101010010",  2265 => b"0000101010001",  2266 => b"0000101010000",  2267 => b"0000101001111",
 2268 => b"0000101001110",  2269 => b"0000101001110",  2270 => b"0000101001101",  2271 => b"0000101001100",
 2272 => b"0000101001011",  2273 => b"0000101001010",  2274 => b"0000101001010",  2275 => b"0000101001001",
 2276 => b"0000101001000",  2277 => b"0000101000111",  2278 => b"0000101000110",  2279 => b"0000101000110",
 2280 => b"0000101000101",  2281 => b"0000101000100",  2282 => b"0000101000011",  2283 => b"0000101000010",
 2284 => b"0000101000010",  2285 => b"0000101000001",  2286 => b"0000101000000",  2287 => b"0000100111111",
 2288 => b"0000100111110",  2289 => b"0000100111110",  2290 => b"0000100111101",  2291 => b"0000100111100",
 2292 => b"0000100111011",  2293 => b"0000100111010",  2294 => b"0000100111010",  2295 => b"0000100111001",
 2296 => b"0000100111000",  2297 => b"0000100110111",  2298 => b"0000100110110",  2299 => b"0000100110110",
 2300 => b"0000100110101",  2301 => b"0000100110100",  2302 => b"0000100110011",  2303 => b"0000100110010",
 2304 => b"0000100110010",  2305 => b"0000100110001",  2306 => b"0000100110000",  2307 => b"0000100101111",
 2308 => b"0000100101110",  2309 => b"0000100101101",  2310 => b"0000100101101",  2311 => b"0000100101100",
 2312 => b"0000100101011",  2313 => b"0000100101010",  2314 => b"0000100101001",  2315 => b"0000100101001",
 2316 => b"0000100101000",  2317 => b"0000100100111",  2318 => b"0000100100110",  2319 => b"0000100100101",
 2320 => b"0000100100101",  2321 => b"0000100100100",  2322 => b"0000100100011",  2323 => b"0000100100010",
 2324 => b"0000100100001",  2325 => b"0000100100001",  2326 => b"0000100100000",  2327 => b"0000100011111",
 2328 => b"0000100011110",  2329 => b"0000100011110",  2330 => b"0000100011101",  2331 => b"0000100011100",
 2332 => b"0000100011011",  2333 => b"0000100011010",  2334 => b"0000100011010",  2335 => b"0000100011001",
 2336 => b"0000100011000",  2337 => b"0000100010111",  2338 => b"0000100010110",  2339 => b"0000100010110",
 2340 => b"0000100010101",  2341 => b"0000100010100",  2342 => b"0000100010011",  2343 => b"0000100010010",
 2344 => b"0000100010010",  2345 => b"0000100010001",  2346 => b"0000100010000",  2347 => b"0000100001111",
 2348 => b"0000100001110",  2349 => b"0000100001110",  2350 => b"0000100001101",  2351 => b"0000100001100",
 2352 => b"0000100001011",  2353 => b"0000100001010",  2354 => b"0000100001010",  2355 => b"0000100001001",
 2356 => b"0000100001000",  2357 => b"0000100000111",  2358 => b"0000100000110",  2359 => b"0000100000110",
 2360 => b"0000100000101",  2361 => b"0000100000100",  2362 => b"0000100000011",  2363 => b"0000100000011",
 2364 => b"0000100000010",  2365 => b"0000100000001",  2366 => b"0000100000000",  2367 => b"0000011111111",
 2368 => b"0000011111111",  2369 => b"0000011111110",  2370 => b"0000011111101",  2371 => b"0000011111100",
 2372 => b"0000011111011",  2373 => b"0000011111011",  2374 => b"0000011111010",  2375 => b"0000011111001",
 2376 => b"0000011111000",  2377 => b"0000011110111",  2378 => b"0000011110111",  2379 => b"0000011110110",
 2380 => b"0000011110101",  2381 => b"0000011110100",  2382 => b"0000011110100",  2383 => b"0000011110011",
 2384 => b"0000011110010",  2385 => b"0000011110001",  2386 => b"0000011110000",  2387 => b"0000011110000",
 2388 => b"0000011101111",  2389 => b"0000011101110",  2390 => b"0000011101101",  2391 => b"0000011101101",
 2392 => b"0000011101100",  2393 => b"0000011101011",  2394 => b"0000011101010",  2395 => b"0000011101001",
 2396 => b"0000011101001",  2397 => b"0000011101000",  2398 => b"0000011100111",  2399 => b"0000011100110",
 2400 => b"0000011100110",  2401 => b"0000011100101",  2402 => b"0000011100100",  2403 => b"0000011100011",
 2404 => b"0000011100010",  2405 => b"0000011100010",  2406 => b"0000011100001",  2407 => b"0000011100000",
 2408 => b"0000011011111",  2409 => b"0000011011111",  2410 => b"0000011011110",  2411 => b"0000011011101",
 2412 => b"0000011011100",  2413 => b"0000011011011",  2414 => b"0000011011011",  2415 => b"0000011011010",
 2416 => b"0000011011001",  2417 => b"0000011011000",  2418 => b"0000011011000",  2419 => b"0000011010111",
 2420 => b"0000011010110",  2421 => b"0000011010101",  2422 => b"0000011010100",  2423 => b"0000011010100",
 2424 => b"0000011010011",  2425 => b"0000011010010",  2426 => b"0000011010001",  2427 => b"0000011010001",
 2428 => b"0000011010000",  2429 => b"0000011001111",  2430 => b"0000011001110",  2431 => b"0000011001110",
 2432 => b"0000011001101",  2433 => b"0000011001100",  2434 => b"0000011001011",  2435 => b"0000011001010",
 2436 => b"0000011001010",  2437 => b"0000011001001",  2438 => b"0000011001000",  2439 => b"0000011000111",
 2440 => b"0000011000111",  2441 => b"0000011000110",  2442 => b"0000011000101",  2443 => b"0000011000100",
 2444 => b"0000011000100",  2445 => b"0000011000011",  2446 => b"0000011000010",  2447 => b"0000011000001",
 2448 => b"0000011000001",  2449 => b"0000011000000",  2450 => b"0000010111111",  2451 => b"0000010111110",
 2452 => b"0000010111110",  2453 => b"0000010111101",  2454 => b"0000010111100",  2455 => b"0000010111011",
 2456 => b"0000010111010",  2457 => b"0000010111010",  2458 => b"0000010111001",  2459 => b"0000010111000",
 2460 => b"0000010110111",  2461 => b"0000010110111",  2462 => b"0000010110110",  2463 => b"0000010110101",
 2464 => b"0000010110100",  2465 => b"0000010110100",  2466 => b"0000010110011",  2467 => b"0000010110010",
 2468 => b"0000010110001",  2469 => b"0000010110001",  2470 => b"0000010110000",  2471 => b"0000010101111",
 2472 => b"0000010101110",  2473 => b"0000010101110",  2474 => b"0000010101101",  2475 => b"0000010101100",
 2476 => b"0000010101011",  2477 => b"0000010101011",  2478 => b"0000010101010",  2479 => b"0000010101001",
 2480 => b"0000010101000",  2481 => b"0000010101000",  2482 => b"0000010100111",  2483 => b"0000010100110",
 2484 => b"0000010100101",  2485 => b"0000010100101",  2486 => b"0000010100100",  2487 => b"0000010100011",
 2488 => b"0000010100010",  2489 => b"0000010100010",  2490 => b"0000010100001",  2491 => b"0000010100000",
 2492 => b"0000010011111",  2493 => b"0000010011111",  2494 => b"0000010011110",  2495 => b"0000010011101",
 2496 => b"0000010011101",  2497 => b"0000010011100",  2498 => b"0000010011011",  2499 => b"0000010011010",
 2500 => b"0000010011010",  2501 => b"0000010011001",  2502 => b"0000010011000",  2503 => b"0000010010111",
 2504 => b"0000010010111",  2505 => b"0000010010110",  2506 => b"0000010010101",  2507 => b"0000010010100",
 2508 => b"0000010010100",  2509 => b"0000010010011",  2510 => b"0000010010010",  2511 => b"0000010010010",
 2512 => b"0000010010001",  2513 => b"0000010010000",  2514 => b"0000010001111",  2515 => b"0000010001111",
 2516 => b"0000010001110",  2517 => b"0000010001101",  2518 => b"0000010001100",  2519 => b"0000010001100",
 2520 => b"0000010001011",  2521 => b"0000010001010",  2522 => b"0000010001001",  2523 => b"0000010001001",
 2524 => b"0000010001000",  2525 => b"0000010000111",  2526 => b"0000010000111",  2527 => b"0000010000110",
 2528 => b"0000010000101",  2529 => b"0000010000100",  2530 => b"0000010000100",  2531 => b"0000010000011",
 2532 => b"0000010000010",  2533 => b"0000010000010",  2534 => b"0000010000001",  2535 => b"0000010000000",
 2536 => b"0000001111111",  2537 => b"0000001111111",  2538 => b"0000001111110",  2539 => b"0000001111101",
 2540 => b"0000001111100",  2541 => b"0000001111100",  2542 => b"0000001111011",  2543 => b"0000001111010",
 2544 => b"0000001111010",  2545 => b"0000001111001",  2546 => b"0000001111000",  2547 => b"0000001110111",
 2548 => b"0000001110111",  2549 => b"0000001110110",  2550 => b"0000001110101",  2551 => b"0000001110101",
 2552 => b"0000001110100",  2553 => b"0000001110011",  2554 => b"0000001110011",  2555 => b"0000001110010",
 2556 => b"0000001110001",  2557 => b"0000001110000",  2558 => b"0000001110000",  2559 => b"0000001101111",
 2560 => b"0000001101110",  2561 => b"0000001101110",  2562 => b"0000001101101",  2563 => b"0000001101100",
 2564 => b"0000001101011",  2565 => b"0000001101011",  2566 => b"0000001101010",  2567 => b"0000001101001",
 2568 => b"0000001101001",  2569 => b"0000001101000",  2570 => b"0000001100111",  2571 => b"0000001100111",
 2572 => b"0000001100110",  2573 => b"0000001100101",  2574 => b"0000001100100",  2575 => b"0000001100100",
 2576 => b"0000001100011",  2577 => b"0000001100010",  2578 => b"0000001100010",  2579 => b"0000001100001",
 2580 => b"0000001100000",  2581 => b"0000001100000",  2582 => b"0000001011111",  2583 => b"0000001011110",
 2584 => b"0000001011110",  2585 => b"0000001011101",  2586 => b"0000001011100",  2587 => b"0000001011011",
 2588 => b"0000001011011",  2589 => b"0000001011010",  2590 => b"0000001011001",  2591 => b"0000001011001",
 2592 => b"0000001011000",  2593 => b"0000001010111",  2594 => b"0000001010111",  2595 => b"0000001010110",
 2596 => b"0000001010101",  2597 => b"0000001010101",  2598 => b"0000001010100",  2599 => b"0000001010011",
 2600 => b"0000001010011",  2601 => b"0000001010010",  2602 => b"0000001010001",  2603 => b"0000001010000",
 2604 => b"0000001010000",  2605 => b"0000001001111",  2606 => b"0000001001110",  2607 => b"0000001001110",
 2608 => b"0000001001101",  2609 => b"0000001001100",  2610 => b"0000001001100",  2611 => b"0000001001011",
 2612 => b"0000001001010",  2613 => b"0000001001010",  2614 => b"0000001001001",  2615 => b"0000001001000",
 2616 => b"0000001001000",  2617 => b"0000001000111",  2618 => b"0000001000110",  2619 => b"0000001000110",
 2620 => b"0000001000101",  2621 => b"0000001000100",  2622 => b"0000001000100",  2623 => b"0000001000011",
 2624 => b"0000001000010",  2625 => b"0000001000010",  2626 => b"0000001000001",  2627 => b"0000001000000",
 2628 => b"0000001000000",  2629 => b"0000000111111",  2630 => b"0000000111110",  2631 => b"0000000111110",
 2632 => b"0000000111101",  2633 => b"0000000111100",  2634 => b"0000000111100",  2635 => b"0000000111011",
 2636 => b"0000000111010",  2637 => b"0000000111010",  2638 => b"0000000111001",  2639 => b"0000000111000",
 2640 => b"0000000111000",  2641 => b"0000000110111",  2642 => b"0000000110110",  2643 => b"0000000110110",
 2644 => b"0000000110101",  2645 => b"0000000110101",  2646 => b"0000000110100",  2647 => b"0000000110011",
 2648 => b"0000000110011",  2649 => b"0000000110010",  2650 => b"0000000110001",  2651 => b"0000000110001",
 2652 => b"0000000110000",  2653 => b"0000000101111",  2654 => b"0000000101111",  2655 => b"0000000101110",
 2656 => b"0000000101101",  2657 => b"0000000101101",  2658 => b"0000000101100",  2659 => b"0000000101011",
 2660 => b"0000000101011",  2661 => b"0000000101010",  2662 => b"0000000101010",  2663 => b"0000000101001",
 2664 => b"0000000101000",  2665 => b"0000000101000",  2666 => b"0000000100111",  2667 => b"0000000100110",
 2668 => b"0000000100110",  2669 => b"0000000100101",  2670 => b"0000000100100",  2671 => b"0000000100100",
 2672 => b"0000000100011",  2673 => b"0000000100011",  2674 => b"0000000100010",  2675 => b"0000000100001",
 2676 => b"0000000100001",  2677 => b"0000000100000",  2678 => b"0000000011111",  2679 => b"0000000011111",
 2680 => b"0000000011110",  2681 => b"0000000011101",  2682 => b"0000000011101",  2683 => b"0000000011100",
 2684 => b"0000000011100",  2685 => b"0000000011011",  2686 => b"0000000011010",  2687 => b"0000000011010",
 2688 => b"0000000011001",  2689 => b"0000000011001",  2690 => b"0000000011000",  2691 => b"0000000010111",
 2692 => b"0000000010111",  2693 => b"0000000010110",  2694 => b"0000000010101",  2695 => b"0000000010101",
 2696 => b"0000000010100",  2697 => b"0000000010100",  2698 => b"0000000010011",  2699 => b"0000000010010",
 2700 => b"0000000010010",  2701 => b"0000000010001",  2702 => b"0000000010001",  2703 => b"0000000010000",
 2704 => b"0000000001111",  2705 => b"0000000001111",  2706 => b"0000000001110",  2707 => b"0000000001101",
 2708 => b"0000000001101",  2709 => b"0000000001100",  2710 => b"0000000001100",  2711 => b"0000000001011",
 2712 => b"0000000001010",  2713 => b"0000000001010",  2714 => b"0000000001001",  2715 => b"0000000001001",
 2716 => b"0000000001000",  2717 => b"0000000000111",  2718 => b"0000000000111",  2719 => b"0000000000110",
 2720 => b"0000000000110",  2721 => b"0000000000101",  2722 => b"0000000000100",  2723 => b"0000000000100",
 2724 => b"0000000000011",  2725 => b"0000000000011",  2726 => b"0000000000010",  2727 => b"0000000000001",
 2728 => b"0000000000001",  2729 => b"0000000000000",  2730 => b"0000000000000",  2731 => b"0000000000000",
 2732 => b"0000000000000",  2733 => b"1111111111111",  2734 => b"1111111111110",  2735 => b"1111111111110",
 2736 => b"1111111111101",  2737 => b"1111111111101",  2738 => b"1111111111100",  2739 => b"1111111111011",
 2740 => b"1111111111011",  2741 => b"1111111111010",  2742 => b"1111111111010",  2743 => b"1111111111001",
 2744 => b"1111111111001",  2745 => b"1111111111000",  2746 => b"1111111110111",  2747 => b"1111111110111",
 2748 => b"1111111110110",  2749 => b"1111111110110",  2750 => b"1111111110101",  2751 => b"1111111110100",
 2752 => b"1111111110100",  2753 => b"1111111110011",  2754 => b"1111111110011",  2755 => b"1111111110010",
 2756 => b"1111111110010",  2757 => b"1111111110001",  2758 => b"1111111110001",  2759 => b"1111111110000",
 2760 => b"1111111101111",  2761 => b"1111111101111",  2762 => b"1111111101110",  2763 => b"1111111101110",
 2764 => b"1111111101101",  2765 => b"1111111101101",  2766 => b"1111111101100",  2767 => b"1111111101011",
 2768 => b"1111111101011",  2769 => b"1111111101010",  2770 => b"1111111101010",  2771 => b"1111111101001",
 2772 => b"1111111101001",  2773 => b"1111111101000",  2774 => b"1111111101000",  2775 => b"1111111100111",
 2776 => b"1111111100110",  2777 => b"1111111100110",  2778 => b"1111111100101",  2779 => b"1111111100101",
 2780 => b"1111111100100",  2781 => b"1111111100100",  2782 => b"1111111100011",  2783 => b"1111111100011",
 2784 => b"1111111100010",  2785 => b"1111111100001",  2786 => b"1111111100001",  2787 => b"1111111100000",
 2788 => b"1111111100000",  2789 => b"1111111011111",  2790 => b"1111111011111",  2791 => b"1111111011110",
 2792 => b"1111111011110",  2793 => b"1111111011101",  2794 => b"1111111011101",  2795 => b"1111111011100",
 2796 => b"1111111011100",  2797 => b"1111111011011",  2798 => b"1111111011010",  2799 => b"1111111011010",
 2800 => b"1111111011001",  2801 => b"1111111011001",  2802 => b"1111111011000",  2803 => b"1111111011000",
 2804 => b"1111111010111",  2805 => b"1111111010111",  2806 => b"1111111010110",  2807 => b"1111111010110",
 2808 => b"1111111010101",  2809 => b"1111111010101",  2810 => b"1111111010100",  2811 => b"1111111010100",
 2812 => b"1111111010011",  2813 => b"1111111010011",  2814 => b"1111111010010",  2815 => b"1111111010010",
 2816 => b"1111111010001",  2817 => b"1111111010000",  2818 => b"1111111010000",  2819 => b"1111111001111",
 2820 => b"1111111001111",  2821 => b"1111111001110",  2822 => b"1111111001110",  2823 => b"1111111001101",
 2824 => b"1111111001101",  2825 => b"1111111001100",  2826 => b"1111111001100",  2827 => b"1111111001011",
 2828 => b"1111111001011",  2829 => b"1111111001010",  2830 => b"1111111001010",  2831 => b"1111111001001",
 2832 => b"1111111001001",  2833 => b"1111111001000",  2834 => b"1111111001000",  2835 => b"1111111000111",
 2836 => b"1111111000111",  2837 => b"1111111000110",  2838 => b"1111111000110",  2839 => b"1111111000101",
 2840 => b"1111111000101",  2841 => b"1111111000100",  2842 => b"1111111000100",  2843 => b"1111111000011",
 2844 => b"1111111000011",  2845 => b"1111111000010",  2846 => b"1111111000010",  2847 => b"1111111000001",
 2848 => b"1111111000001",  2849 => b"1111111000000",  2850 => b"1111111000000",  2851 => b"1111110111111",
 2852 => b"1111110111111",  2853 => b"1111110111110",  2854 => b"1111110111110",  2855 => b"1111110111101",
 2856 => b"1111110111101",  2857 => b"1111110111100",  2858 => b"1111110111100",  2859 => b"1111110111100",
 2860 => b"1111110111011",  2861 => b"1111110111011",  2862 => b"1111110111010",  2863 => b"1111110111010",
 2864 => b"1111110111001",  2865 => b"1111110111001",  2866 => b"1111110111000",  2867 => b"1111110111000",
 2868 => b"1111110110111",  2869 => b"1111110110111",  2870 => b"1111110110110",  2871 => b"1111110110110",
 2872 => b"1111110110101",  2873 => b"1111110110101",  2874 => b"1111110110100",  2875 => b"1111110110100",
 2876 => b"1111110110011",  2877 => b"1111110110011",  2878 => b"1111110110011",  2879 => b"1111110110010",
 2880 => b"1111110110010",  2881 => b"1111110110001",  2882 => b"1111110110001",  2883 => b"1111110110000",
 2884 => b"1111110110000",  2885 => b"1111110101111",  2886 => b"1111110101111",  2887 => b"1111110101110",
 2888 => b"1111110101110",  2889 => b"1111110101110",  2890 => b"1111110101101",  2891 => b"1111110101101",
 2892 => b"1111110101100",  2893 => b"1111110101100",  2894 => b"1111110101011",  2895 => b"1111110101011",
 2896 => b"1111110101010",  2897 => b"1111110101010",  2898 => b"1111110101001",  2899 => b"1111110101001",
 2900 => b"1111110101001",  2901 => b"1111110101000",  2902 => b"1111110101000",  2903 => b"1111110100111",
 2904 => b"1111110100111",  2905 => b"1111110100110",  2906 => b"1111110100110",  2907 => b"1111110100101",
 2908 => b"1111110100101",  2909 => b"1111110100101",  2910 => b"1111110100100",  2911 => b"1111110100100",
 2912 => b"1111110100011",  2913 => b"1111110100011",  2914 => b"1111110100010",  2915 => b"1111110100010",
 2916 => b"1111110100010",  2917 => b"1111110100001",  2918 => b"1111110100001",  2919 => b"1111110100000",
 2920 => b"1111110100000",  2921 => b"1111110011111",  2922 => b"1111110011111",  2923 => b"1111110011111",
 2924 => b"1111110011110",  2925 => b"1111110011110",  2926 => b"1111110011101",  2927 => b"1111110011101",
 2928 => b"1111110011101",  2929 => b"1111110011100",  2930 => b"1111110011100",  2931 => b"1111110011011",
 2932 => b"1111110011011",  2933 => b"1111110011010",  2934 => b"1111110011010",  2935 => b"1111110011010",
 2936 => b"1111110011001",  2937 => b"1111110011001",  2938 => b"1111110011000",  2939 => b"1111110011000",
 2940 => b"1111110011000",  2941 => b"1111110010111",  2942 => b"1111110010111",  2943 => b"1111110010110",
 2944 => b"1111110010110",  2945 => b"1111110010110",  2946 => b"1111110010101",  2947 => b"1111110010101",
 2948 => b"1111110010100",  2949 => b"1111110010100",  2950 => b"1111110010100",  2951 => b"1111110010011",
 2952 => b"1111110010011",  2953 => b"1111110010010",  2954 => b"1111110010010",  2955 => b"1111110010010",
 2956 => b"1111110010001",  2957 => b"1111110010001",  2958 => b"1111110010000",  2959 => b"1111110010000",
 2960 => b"1111110010000",  2961 => b"1111110001111",  2962 => b"1111110001111",  2963 => b"1111110001111",
 2964 => b"1111110001110",  2965 => b"1111110001110",  2966 => b"1111110001101",  2967 => b"1111110001101",
 2968 => b"1111110001101",  2969 => b"1111110001100",  2970 => b"1111110001100",  2971 => b"1111110001011",
 2972 => b"1111110001011",  2973 => b"1111110001011",  2974 => b"1111110001010",  2975 => b"1111110001010",
 2976 => b"1111110001010",  2977 => b"1111110001001",  2978 => b"1111110001001",  2979 => b"1111110001000",
 2980 => b"1111110001000",  2981 => b"1111110001000",  2982 => b"1111110000111",  2983 => b"1111110000111",
 2984 => b"1111110000111",  2985 => b"1111110000110",  2986 => b"1111110000110",  2987 => b"1111110000110",
 2988 => b"1111110000101",  2989 => b"1111110000101",  2990 => b"1111110000100",  2991 => b"1111110000100",
 2992 => b"1111110000100",  2993 => b"1111110000011",  2994 => b"1111110000011",  2995 => b"1111110000011",
 2996 => b"1111110000010",  2997 => b"1111110000010",  2998 => b"1111110000010",  2999 => b"1111110000001",
 3000 => b"1111110000001",  3001 => b"1111110000001",  3002 => b"1111110000000",  3003 => b"1111110000000",
 3004 => b"1111110000000",  3005 => b"1111101111111",  3006 => b"1111101111111",  3007 => b"1111101111111",
 3008 => b"1111101111110",  3009 => b"1111101111110",  3010 => b"1111101111110",  3011 => b"1111101111101",
 3012 => b"1111101111101",  3013 => b"1111101111101",  3014 => b"1111101111100",  3015 => b"1111101111100",
 3016 => b"1111101111100",  3017 => b"1111101111011",  3018 => b"1111101111011",  3019 => b"1111101111011",
 3020 => b"1111101111010",  3021 => b"1111101111010",  3022 => b"1111101111010",  3023 => b"1111101111001",
 3024 => b"1111101111001",  3025 => b"1111101111001",  3026 => b"1111101111000",  3027 => b"1111101111000",
 3028 => b"1111101111000",  3029 => b"1111101110111",  3030 => b"1111101110111",  3031 => b"1111101110111",
 3032 => b"1111101110110",  3033 => b"1111101110110",  3034 => b"1111101110110",  3035 => b"1111101110101",
 3036 => b"1111101110101",  3037 => b"1111101110101",  3038 => b"1111101110100",  3039 => b"1111101110100",
 3040 => b"1111101110100",  3041 => b"1111101110100",  3042 => b"1111101110011",  3043 => b"1111101110011",
 3044 => b"1111101110011",  3045 => b"1111101110010",  3046 => b"1111101110010",  3047 => b"1111101110010",
 3048 => b"1111101110001",  3049 => b"1111101110001",  3050 => b"1111101110001",  3051 => b"1111101110000",
 3052 => b"1111101110000",  3053 => b"1111101110000",  3054 => b"1111101110000",  3055 => b"1111101101111",
 3056 => b"1111101101111",  3057 => b"1111101101111",  3058 => b"1111101101110",  3059 => b"1111101101110",
 3060 => b"1111101101110",  3061 => b"1111101101110",  3062 => b"1111101101101",  3063 => b"1111101101101",
 3064 => b"1111101101101",  3065 => b"1111101101100",  3066 => b"1111101101100",  3067 => b"1111101101100",
 3068 => b"1111101101100",  3069 => b"1111101101011",  3070 => b"1111101101011",  3071 => b"1111101101011",
 3072 => b"1111101101010",  3073 => b"1111101101010",  3074 => b"1111101101010",  3075 => b"1111101101010",
 3076 => b"1111101101001",  3077 => b"1111101101001",  3078 => b"1111101101001",  3079 => b"1111101101001",
 3080 => b"1111101101000",  3081 => b"1111101101000",  3082 => b"1111101101000",  3083 => b"1111101100111",
 3084 => b"1111101100111",  3085 => b"1111101100111",  3086 => b"1111101100111",  3087 => b"1111101100110",
 3088 => b"1111101100110",  3089 => b"1111101100110",  3090 => b"1111101100110",  3091 => b"1111101100101",
 3092 => b"1111101100101",  3093 => b"1111101100101",  3094 => b"1111101100101",  3095 => b"1111101100100",
 3096 => b"1111101100100",  3097 => b"1111101100100",  3098 => b"1111101100100",  3099 => b"1111101100011",
 3100 => b"1111101100011",  3101 => b"1111101100011",  3102 => b"1111101100011",  3103 => b"1111101100010",
 3104 => b"1111101100010",  3105 => b"1111101100010",  3106 => b"1111101100010",  3107 => b"1111101100001",
 3108 => b"1111101100001",  3109 => b"1111101100001",  3110 => b"1111101100001",  3111 => b"1111101100000",
 3112 => b"1111101100000",  3113 => b"1111101100000",  3114 => b"1111101100000",  3115 => b"1111101011111",
 3116 => b"1111101011111",  3117 => b"1111101011111",  3118 => b"1111101011111",  3119 => b"1111101011110",
 3120 => b"1111101011110",  3121 => b"1111101011110",  3122 => b"1111101011110",  3123 => b"1111101011110",
 3124 => b"1111101011101",  3125 => b"1111101011101",  3126 => b"1111101011101",  3127 => b"1111101011101",
 3128 => b"1111101011100",  3129 => b"1111101011100",  3130 => b"1111101011100",  3131 => b"1111101011100",
 3132 => b"1111101011100",  3133 => b"1111101011011",  3134 => b"1111101011011",  3135 => b"1111101011011",
 3136 => b"1111101011011",  3137 => b"1111101011011",  3138 => b"1111101011010",  3139 => b"1111101011010",
 3140 => b"1111101011010",  3141 => b"1111101011010",  3142 => b"1111101011001",  3143 => b"1111101011001",
 3144 => b"1111101011001",  3145 => b"1111101011001",  3146 => b"1111101011001",  3147 => b"1111101011000",
 3148 => b"1111101011000",  3149 => b"1111101011000",  3150 => b"1111101011000",  3151 => b"1111101011000",
 3152 => b"1111101010111",  3153 => b"1111101010111",  3154 => b"1111101010111",  3155 => b"1111101010111",
 3156 => b"1111101010111",  3157 => b"1111101010110",  3158 => b"1111101010110",  3159 => b"1111101010110",
 3160 => b"1111101010110",  3161 => b"1111101010110",  3162 => b"1111101010110",  3163 => b"1111101010101",
 3164 => b"1111101010101",  3165 => b"1111101010101",  3166 => b"1111101010101",  3167 => b"1111101010101",
 3168 => b"1111101010100",  3169 => b"1111101010100",  3170 => b"1111101010100",  3171 => b"1111101010100",
 3172 => b"1111101010100",  3173 => b"1111101010011",  3174 => b"1111101010011",  3175 => b"1111101010011",
 3176 => b"1111101010011",  3177 => b"1111101010011",  3178 => b"1111101010011",  3179 => b"1111101010010",
 3180 => b"1111101010010",  3181 => b"1111101010010",  3182 => b"1111101010010",  3183 => b"1111101010010",
 3184 => b"1111101010010",  3185 => b"1111101010001",  3186 => b"1111101010001",  3187 => b"1111101010001",
 3188 => b"1111101010001",  3189 => b"1111101010001",  3190 => b"1111101010001",  3191 => b"1111101010000",
 3192 => b"1111101010000",  3193 => b"1111101010000",  3194 => b"1111101010000",  3195 => b"1111101010000",
 3196 => b"1111101010000",  3197 => b"1111101010000",  3198 => b"1111101001111",  3199 => b"1111101001111",
 3200 => b"1111101001111",  3201 => b"1111101001111",  3202 => b"1111101001111",  3203 => b"1111101001111",
 3204 => b"1111101001110",  3205 => b"1111101001110",  3206 => b"1111101001110",  3207 => b"1111101001110",
 3208 => b"1111101001110",  3209 => b"1111101001110",  3210 => b"1111101001110",  3211 => b"1111101001101",
 3212 => b"1111101001101",  3213 => b"1111101001101",  3214 => b"1111101001101",  3215 => b"1111101001101",
 3216 => b"1111101001101",  3217 => b"1111101001101",  3218 => b"1111101001101",  3219 => b"1111101001100",
 3220 => b"1111101001100",  3221 => b"1111101001100",  3222 => b"1111101001100",  3223 => b"1111101001100",
 3224 => b"1111101001100",  3225 => b"1111101001100",  3226 => b"1111101001100",  3227 => b"1111101001011",
 3228 => b"1111101001011",  3229 => b"1111101001011",  3230 => b"1111101001011",  3231 => b"1111101001011",
 3232 => b"1111101001011",  3233 => b"1111101001011",  3234 => b"1111101001011",  3235 => b"1111101001010",
 3236 => b"1111101001010",  3237 => b"1111101001010",  3238 => b"1111101001010",  3239 => b"1111101001010",
 3240 => b"1111101001010",  3241 => b"1111101001010",  3242 => b"1111101001010",  3243 => b"1111101001010",
 3244 => b"1111101001001",  3245 => b"1111101001001",  3246 => b"1111101001001",  3247 => b"1111101001001",
 3248 => b"1111101001001",  3249 => b"1111101001001",  3250 => b"1111101001001",  3251 => b"1111101001001",
 3252 => b"1111101001001",  3253 => b"1111101001001",  3254 => b"1111101001000",  3255 => b"1111101001000",
 3256 => b"1111101001000",  3257 => b"1111101001000",  3258 => b"1111101001000",  3259 => b"1111101001000",
 3260 => b"1111101001000",  3261 => b"1111101001000",  3262 => b"1111101001000",  3263 => b"1111101001000",
 3264 => b"1111101001000",  3265 => b"1111101000111",  3266 => b"1111101000111",  3267 => b"1111101000111",
 3268 => b"1111101000111",  3269 => b"1111101000111",  3270 => b"1111101000111",  3271 => b"1111101000111",
 3272 => b"1111101000111",  3273 => b"1111101000111",  3274 => b"1111101000111",  3275 => b"1111101000111",
 3276 => b"1111101000111",  3277 => b"1111101000110",  3278 => b"1111101000110",  3279 => b"1111101000110",
 3280 => b"1111101000110",  3281 => b"1111101000110",  3282 => b"1111101000110",  3283 => b"1111101000110",
 3284 => b"1111101000110",  3285 => b"1111101000110",  3286 => b"1111101000110",  3287 => b"1111101000110",
 3288 => b"1111101000110",  3289 => b"1111101000110",  3290 => b"1111101000110",  3291 => b"1111101000110",
 3292 => b"1111101000101",  3293 => b"1111101000101",  3294 => b"1111101000101",  3295 => b"1111101000101",
 3296 => b"1111101000101",  3297 => b"1111101000101",  3298 => b"1111101000101",  3299 => b"1111101000101",
 3300 => b"1111101000101",  3301 => b"1111101000101",  3302 => b"1111101000101",  3303 => b"1111101000101",
 3304 => b"1111101000101",  3305 => b"1111101000101",  3306 => b"1111101000101",  3307 => b"1111101000101",
 3308 => b"1111101000101",  3309 => b"1111101000101",  3310 => b"1111101000101",  3311 => b"1111101000100",
 3312 => b"1111101000100",  3313 => b"1111101000100",  3314 => b"1111101000100",  3315 => b"1111101000100",
 3316 => b"1111101000100",  3317 => b"1111101000100",  3318 => b"1111101000100",  3319 => b"1111101000100",
 3320 => b"1111101000100",  3321 => b"1111101000100",  3322 => b"1111101000100",  3323 => b"1111101000100",
 3324 => b"1111101000100",  3325 => b"1111101000100",  3326 => b"1111101000100",  3327 => b"1111101000100",
 3328 => b"1111101000100",  3329 => b"1111101000100",  3330 => b"1111101000100",  3331 => b"1111101000100",
 3332 => b"1111101000100",  3333 => b"1111101000100",  3334 => b"1111101000100",  3335 => b"1111101000100",
 3336 => b"1111101000100",  3337 => b"1111101000100",  3338 => b"1111101000100",  3339 => b"1111101000100",
 3340 => b"1111101000100",  3341 => b"1111101000100",  3342 => b"1111101000100",  3343 => b"1111101000100",
 3344 => b"1111101000100",  3345 => b"1111101000100",  3346 => b"1111101000100",  3347 => b"1111101000100",
 3348 => b"1111101000100",  3349 => b"1111101000100",  3350 => b"1111101000100",  3351 => b"1111101000100",
 3352 => b"1111101000100",  3353 => b"1111101000100",  3354 => b"1111101000100",  3355 => b"1111101000100",
 3356 => b"1111101000100",  3357 => b"1111101000100",  3358 => b"1111101000100",  3359 => b"1111101000100",
 3360 => b"1111101000100",  3361 => b"1111101000100",  3362 => b"1111101000100",  3363 => b"1111101000100",
 3364 => b"1111101000100",  3365 => b"1111101000100",  3366 => b"1111101000100",  3367 => b"1111101000100",
 3368 => b"1111101000100",  3369 => b"1111101000100",  3370 => b"1111101000100",  3371 => b"1111101000100",
 3372 => b"1111101000100",  3373 => b"1111101000100",  3374 => b"1111101000100",  3375 => b"1111101000100",
 3376 => b"1111101000100",  3377 => b"1111101000100",  3378 => b"1111101000100",  3379 => b"1111101000100",
 3380 => b"1111101000100",  3381 => b"1111101000100",  3382 => b"1111101000100",  3383 => b"1111101000100",
 3384 => b"1111101000100",  3385 => b"1111101000100",  3386 => b"1111101000100",  3387 => b"1111101000100",
 3388 => b"1111101000100",  3389 => b"1111101000100",  3390 => b"1111101000100",  3391 => b"1111101000100",
 3392 => b"1111101000100",  3393 => b"1111101000100",  3394 => b"1111101000100",  3395 => b"1111101000100",
 3396 => b"1111101000100",  3397 => b"1111101000100",  3398 => b"1111101000100",  3399 => b"1111101000100",
 3400 => b"1111101000100",  3401 => b"1111101000101",  3402 => b"1111101000101",  3403 => b"1111101000101",
 3404 => b"1111101000101",  3405 => b"1111101000101",  3406 => b"1111101000101",  3407 => b"1111101000101",
 3408 => b"1111101000101",  3409 => b"1111101000101",  3410 => b"1111101000101",  3411 => b"1111101000101",
 3412 => b"1111101000101",  3413 => b"1111101000101",  3414 => b"1111101000101",  3415 => b"1111101000101",
 3416 => b"1111101000101",  3417 => b"1111101000101",  3418 => b"1111101000101",  3419 => b"1111101000101",
 3420 => b"1111101000101",  3421 => b"1111101000110",  3422 => b"1111101000110",  3423 => b"1111101000110",
 3424 => b"1111101000110",  3425 => b"1111101000110",  3426 => b"1111101000110",  3427 => b"1111101000110",
 3428 => b"1111101000110",  3429 => b"1111101000110",  3430 => b"1111101000110",  3431 => b"1111101000110",
 3432 => b"1111101000110",  3433 => b"1111101000110",  3434 => b"1111101000110",  3435 => b"1111101000110",
 3436 => b"1111101000111",  3437 => b"1111101000111",  3438 => b"1111101000111",  3439 => b"1111101000111",
 3440 => b"1111101000111",  3441 => b"1111101000111",  3442 => b"1111101000111",  3443 => b"1111101000111",
 3444 => b"1111101000111",  3445 => b"1111101000111",  3446 => b"1111101000111",  3447 => b"1111101000111",
 3448 => b"1111101000111",  3449 => b"1111101001000",  3450 => b"1111101001000",  3451 => b"1111101001000",
 3452 => b"1111101001000",  3453 => b"1111101001000",  3454 => b"1111101001000",  3455 => b"1111101001000",
 3456 => b"1111101001000",  3457 => b"1111101001000",  3458 => b"1111101001000",  3459 => b"1111101001000",
 3460 => b"1111101001001",  3461 => b"1111101001001",  3462 => b"1111101001001",  3463 => b"1111101001001",
 3464 => b"1111101001001",  3465 => b"1111101001001",  3466 => b"1111101001001",  3467 => b"1111101001001",
 3468 => b"1111101001001",  3469 => b"1111101001001",  3470 => b"1111101001010",  3471 => b"1111101001010",
 3472 => b"1111101001010",  3473 => b"1111101001010",  3474 => b"1111101001010",  3475 => b"1111101001010",
 3476 => b"1111101001010",  3477 => b"1111101001010",  3478 => b"1111101001010",  3479 => b"1111101001010",
 3480 => b"1111101001011",  3481 => b"1111101001011",  3482 => b"1111101001011",  3483 => b"1111101001011",
 3484 => b"1111101001011",  3485 => b"1111101001011",  3486 => b"1111101001011",  3487 => b"1111101001011",
 3488 => b"1111101001100",  3489 => b"1111101001100",  3490 => b"1111101001100",  3491 => b"1111101001100",
 3492 => b"1111101001100",  3493 => b"1111101001100",  3494 => b"1111101001100",  3495 => b"1111101001100",
 3496 => b"1111101001100",  3497 => b"1111101001101",  3498 => b"1111101001101",  3499 => b"1111101001101",
 3500 => b"1111101001101",  3501 => b"1111101001101",  3502 => b"1111101001101",  3503 => b"1111101001101",
 3504 => b"1111101001101",  3505 => b"1111101001110",  3506 => b"1111101001110",  3507 => b"1111101001110",
 3508 => b"1111101001110",  3509 => b"1111101001110",  3510 => b"1111101001110",  3511 => b"1111101001110",
 3512 => b"1111101001111",  3513 => b"1111101001111",  3514 => b"1111101001111",  3515 => b"1111101001111",
 3516 => b"1111101001111",  3517 => b"1111101001111",  3518 => b"1111101001111",  3519 => b"1111101010000",
 3520 => b"1111101010000",  3521 => b"1111101010000",  3522 => b"1111101010000",  3523 => b"1111101010000",
 3524 => b"1111101010000",  3525 => b"1111101010000",  3526 => b"1111101010001",  3527 => b"1111101010001",
 3528 => b"1111101010001",  3529 => b"1111101010001",  3530 => b"1111101010001",  3531 => b"1111101010001",
 3532 => b"1111101010001",  3533 => b"1111101010010",  3534 => b"1111101010010",  3535 => b"1111101010010",
 3536 => b"1111101010010",  3537 => b"1111101010010",  3538 => b"1111101010010",  3539 => b"1111101010011",
 3540 => b"1111101010011",  3541 => b"1111101010011",  3542 => b"1111101010011",  3543 => b"1111101010011",
 3544 => b"1111101010011",  3545 => b"1111101010100",  3546 => b"1111101010100",  3547 => b"1111101010100",
 3548 => b"1111101010100",  3549 => b"1111101010100",  3550 => b"1111101010100",  3551 => b"1111101010101",
 3552 => b"1111101010101",  3553 => b"1111101010101",  3554 => b"1111101010101",  3555 => b"1111101010101",
 3556 => b"1111101010101",  3557 => b"1111101010110",  3558 => b"1111101010110",  3559 => b"1111101010110",
 3560 => b"1111101010110",  3561 => b"1111101010110",  3562 => b"1111101010110",  3563 => b"1111101010111",
 3564 => b"1111101010111",  3565 => b"1111101010111",  3566 => b"1111101010111",  3567 => b"1111101010111",
 3568 => b"1111101010111",  3569 => b"1111101011000",  3570 => b"1111101011000",  3571 => b"1111101011000",
 3572 => b"1111101011000",  3573 => b"1111101011000",  3574 => b"1111101011001",  3575 => b"1111101011001",
 3576 => b"1111101011001",  3577 => b"1111101011001",  3578 => b"1111101011001",  3579 => b"1111101011010",
 3580 => b"1111101011010",  3581 => b"1111101011010",  3582 => b"1111101011010",  3583 => b"1111101011010",
 3584 => b"1111101011010",  3585 => b"1111101011011",  3586 => b"1111101011011",  3587 => b"1111101011011",
 3588 => b"1111101011011",  3589 => b"1111101011011",  3590 => b"1111101011100",  3591 => b"1111101011100",
 3592 => b"1111101011100",  3593 => b"1111101011100",  3594 => b"1111101011100",  3595 => b"1111101011101",
 3596 => b"1111101011101",  3597 => b"1111101011101",  3598 => b"1111101011101",  3599 => b"1111101011101",
 3600 => b"1111101011110",  3601 => b"1111101011110",  3602 => b"1111101011110",  3603 => b"1111101011110",
 3604 => b"1111101011110",  3605 => b"1111101011111",  3606 => b"1111101011111",  3607 => b"1111101011111",
 3608 => b"1111101011111",  3609 => b"1111101100000",  3610 => b"1111101100000",  3611 => b"1111101100000",
 3612 => b"1111101100000",  3613 => b"1111101100000",  3614 => b"1111101100001",  3615 => b"1111101100001",
 3616 => b"1111101100001",  3617 => b"1111101100001",  3618 => b"1111101100001",  3619 => b"1111101100010",
 3620 => b"1111101100010",  3621 => b"1111101100010",  3622 => b"1111101100010",  3623 => b"1111101100011",
 3624 => b"1111101100011",  3625 => b"1111101100011",  3626 => b"1111101100011",  3627 => b"1111101100011",
 3628 => b"1111101100100",  3629 => b"1111101100100",  3630 => b"1111101100100",  3631 => b"1111101100100",
 3632 => b"1111101100101",  3633 => b"1111101100101",  3634 => b"1111101100101",  3635 => b"1111101100101",
 3636 => b"1111101100101",  3637 => b"1111101100110",  3638 => b"1111101100110",  3639 => b"1111101100110",
 3640 => b"1111101100110",  3641 => b"1111101100111",  3642 => b"1111101100111",  3643 => b"1111101100111",
 3644 => b"1111101100111",  3645 => b"1111101101000",  3646 => b"1111101101000",  3647 => b"1111101101000",
 3648 => b"1111101101000",  3649 => b"1111101101001",  3650 => b"1111101101001",  3651 => b"1111101101001",
 3652 => b"1111101101001",  3653 => b"1111101101001",  3654 => b"1111101101010",  3655 => b"1111101101010",
 3656 => b"1111101101010",  3657 => b"1111101101010",  3658 => b"1111101101011",  3659 => b"1111101101011",
 3660 => b"1111101101011",  3661 => b"1111101101011",  3662 => b"1111101101100",  3663 => b"1111101101100",
 3664 => b"1111101101100",  3665 => b"1111101101100",  3666 => b"1111101101101",  3667 => b"1111101101101",
 3668 => b"1111101101101",  3669 => b"1111101101101",  3670 => b"1111101101110",  3671 => b"1111101101110",
 3672 => b"1111101101110",  3673 => b"1111101101110",  3674 => b"1111101101111",  3675 => b"1111101101111",
 3676 => b"1111101101111",  3677 => b"1111101101111",  3678 => b"1111101110000",  3679 => b"1111101110000",
 3680 => b"1111101110000",  3681 => b"1111101110000",  3682 => b"1111101110001",  3683 => b"1111101110001",
 3684 => b"1111101110001",  3685 => b"1111101110010",  3686 => b"1111101110010",  3687 => b"1111101110010",
 3688 => b"1111101110010",  3689 => b"1111101110011",  3690 => b"1111101110011",  3691 => b"1111101110011",
 3692 => b"1111101110011",  3693 => b"1111101110100",  3694 => b"1111101110100",  3695 => b"1111101110100",
 3696 => b"1111101110100",  3697 => b"1111101110101",  3698 => b"1111101110101",  3699 => b"1111101110101",
 3700 => b"1111101110110",  3701 => b"1111101110110",  3702 => b"1111101110110",  3703 => b"1111101110110",
 3704 => b"1111101110111",  3705 => b"1111101110111",  3706 => b"1111101110111",  3707 => b"1111101110111",
 3708 => b"1111101111000",  3709 => b"1111101111000",  3710 => b"1111101111000",  3711 => b"1111101111001",
 3712 => b"1111101111001",  3713 => b"1111101111001",  3714 => b"1111101111001",  3715 => b"1111101111010",
 3716 => b"1111101111010",  3717 => b"1111101111010",  3718 => b"1111101111010",  3719 => b"1111101111011",
 3720 => b"1111101111011",  3721 => b"1111101111011",  3722 => b"1111101111100",  3723 => b"1111101111100",
 3724 => b"1111101111100",  3725 => b"1111101111100",  3726 => b"1111101111101",  3727 => b"1111101111101",
 3728 => b"1111101111101",  3729 => b"1111101111110",  3730 => b"1111101111110",  3731 => b"1111101111110",
 3732 => b"1111101111110",  3733 => b"1111101111111",  3734 => b"1111101111111",  3735 => b"1111101111111",
 3736 => b"1111110000000",  3737 => b"1111110000000",  3738 => b"1111110000000",  3739 => b"1111110000001",
 3740 => b"1111110000001",  3741 => b"1111110000001",  3742 => b"1111110000001",  3743 => b"1111110000010",
 3744 => b"1111110000010",  3745 => b"1111110000010",  3746 => b"1111110000011",  3747 => b"1111110000011",
 3748 => b"1111110000011",  3749 => b"1111110000011",  3750 => b"1111110000100",  3751 => b"1111110000100",
 3752 => b"1111110000100",  3753 => b"1111110000101",  3754 => b"1111110000101",  3755 => b"1111110000101",
 3756 => b"1111110000110",  3757 => b"1111110000110",  3758 => b"1111110000110",  3759 => b"1111110000110",
 3760 => b"1111110000111",  3761 => b"1111110000111",  3762 => b"1111110000111",  3763 => b"1111110001000",
 3764 => b"1111110001000",  3765 => b"1111110001000",  3766 => b"1111110001001",  3767 => b"1111110001001",
 3768 => b"1111110001001",  3769 => b"1111110001010",  3770 => b"1111110001010",  3771 => b"1111110001010",
 3772 => b"1111110001010",  3773 => b"1111110001011",  3774 => b"1111110001011",  3775 => b"1111110001011",
 3776 => b"1111110001100",  3777 => b"1111110001100",  3778 => b"1111110001100",  3779 => b"1111110001101",
 3780 => b"1111110001101",  3781 => b"1111110001101",  3782 => b"1111110001110",  3783 => b"1111110001110",
 3784 => b"1111110001110",  3785 => b"1111110001111",  3786 => b"1111110001111",  3787 => b"1111110001111",
 3788 => b"1111110001111",  3789 => b"1111110010000",  3790 => b"1111110010000",  3791 => b"1111110010000",
 3792 => b"1111110010001",  3793 => b"1111110010001",  3794 => b"1111110010001",  3795 => b"1111110010010",
 3796 => b"1111110010010",  3797 => b"1111110010010",  3798 => b"1111110010011",  3799 => b"1111110010011",
 3800 => b"1111110010011",  3801 => b"1111110010100",  3802 => b"1111110010100",  3803 => b"1111110010100",
 3804 => b"1111110010101",  3805 => b"1111110010101",  3806 => b"1111110010101",  3807 => b"1111110010110",
 3808 => b"1111110010110",  3809 => b"1111110010110",  3810 => b"1111110010111",  3811 => b"1111110010111",
 3812 => b"1111110010111",  3813 => b"1111110011000",  3814 => b"1111110011000",  3815 => b"1111110011000",
 3816 => b"1111110011001",  3817 => b"1111110011001",  3818 => b"1111110011001",  3819 => b"1111110011010",
 3820 => b"1111110011010",  3821 => b"1111110011010",  3822 => b"1111110011011",  3823 => b"1111110011011",
 3824 => b"1111110011011",  3825 => b"1111110011100",  3826 => b"1111110011100",  3827 => b"1111110011100",
 3828 => b"1111110011101",  3829 => b"1111110011101",  3830 => b"1111110011101",  3831 => b"1111110011110",
 3832 => b"1111110011110",  3833 => b"1111110011110",  3834 => b"1111110011111",  3835 => b"1111110011111",
 3836 => b"1111110011111",  3837 => b"1111110100000",  3838 => b"1111110100000",  3839 => b"1111110100000",
 3840 => b"1111110100001",  3841 => b"1111110100001",  3842 => b"1111110100001",  3843 => b"1111110100010",
 3844 => b"1111110100010",  3845 => b"1111110100010",  3846 => b"1111110100011",  3847 => b"1111110100011",
 3848 => b"1111110100011",  3849 => b"1111110100100",  3850 => b"1111110100100",  3851 => b"1111110100100",
 3852 => b"1111110100101",  3853 => b"1111110100101",  3854 => b"1111110100101",  3855 => b"1111110100110",
 3856 => b"1111110100110",  3857 => b"1111110100110",  3858 => b"1111110100111",  3859 => b"1111110100111",
 3860 => b"1111110101000",  3861 => b"1111110101000",  3862 => b"1111110101000",  3863 => b"1111110101001",
 3864 => b"1111110101001",  3865 => b"1111110101001",  3866 => b"1111110101010",  3867 => b"1111110101010",
 3868 => b"1111110101010",  3869 => b"1111110101011",  3870 => b"1111110101011",  3871 => b"1111110101011",
 3872 => b"1111110101100",  3873 => b"1111110101100",  3874 => b"1111110101100",  3875 => b"1111110101101",
 3876 => b"1111110101101",  3877 => b"1111110101101",  3878 => b"1111110101110",  3879 => b"1111110101110",
 3880 => b"1111110101111",  3881 => b"1111110101111",  3882 => b"1111110101111",  3883 => b"1111110110000",
 3884 => b"1111110110000",  3885 => b"1111110110000",  3886 => b"1111110110001",  3887 => b"1111110110001",
 3888 => b"1111110110001",  3889 => b"1111110110010",  3890 => b"1111110110010",  3891 => b"1111110110010",
 3892 => b"1111110110011",  3893 => b"1111110110011",  3894 => b"1111110110100",  3895 => b"1111110110100",
 3896 => b"1111110110100",  3897 => b"1111110110101",  3898 => b"1111110110101",  3899 => b"1111110110101",
 3900 => b"1111110110110",  3901 => b"1111110110110",  3902 => b"1111110110110",  3903 => b"1111110110111",
 3904 => b"1111110110111",  3905 => b"1111110111000",  3906 => b"1111110111000",  3907 => b"1111110111000",
 3908 => b"1111110111001",  3909 => b"1111110111001",  3910 => b"1111110111001",  3911 => b"1111110111010",
 3912 => b"1111110111010",  3913 => b"1111110111010",  3914 => b"1111110111011",  3915 => b"1111110111011",
 3916 => b"1111110111100",  3917 => b"1111110111100",  3918 => b"1111110111100",  3919 => b"1111110111101",
 3920 => b"1111110111101",  3921 => b"1111110111101",  3922 => b"1111110111110",  3923 => b"1111110111110",
 3924 => b"1111110111110",  3925 => b"1111110111111",  3926 => b"1111110111111",  3927 => b"1111111000000",
 3928 => b"1111111000000",  3929 => b"1111111000000",  3930 => b"1111111000001",  3931 => b"1111111000001",
 3932 => b"1111111000001",  3933 => b"1111111000010",  3934 => b"1111111000010",  3935 => b"1111111000011",
 3936 => b"1111111000011",  3937 => b"1111111000011",  3938 => b"1111111000100",  3939 => b"1111111000100",
 3940 => b"1111111000100",  3941 => b"1111111000101",  3942 => b"1111111000101",  3943 => b"1111111000110",
 3944 => b"1111111000110",  3945 => b"1111111000110",  3946 => b"1111111000111",  3947 => b"1111111000111",
 3948 => b"1111111000111",  3949 => b"1111111001000",  3950 => b"1111111001000",  3951 => b"1111111001001",
 3952 => b"1111111001001",  3953 => b"1111111001001",  3954 => b"1111111001010",  3955 => b"1111111001010",
 3956 => b"1111111001010",  3957 => b"1111111001011",  3958 => b"1111111001011",  3959 => b"1111111001100",
 3960 => b"1111111001100",  3961 => b"1111111001100",  3962 => b"1111111001101",  3963 => b"1111111001101",
 3964 => b"1111111001101",  3965 => b"1111111001110",  3966 => b"1111111001110",  3967 => b"1111111001111",
 3968 => b"1111111001111",  3969 => b"1111111001111",  3970 => b"1111111010000",  3971 => b"1111111010000",
 3972 => b"1111111010001",  3973 => b"1111111010001",  3974 => b"1111111010001",  3975 => b"1111111010010",
 3976 => b"1111111010010",  3977 => b"1111111010010",  3978 => b"1111111010011",  3979 => b"1111111010011",
 3980 => b"1111111010100",  3981 => b"1111111010100",  3982 => b"1111111010100",  3983 => b"1111111010101",
 3984 => b"1111111010101",  3985 => b"1111111010101",  3986 => b"1111111010110",  3987 => b"1111111010110",
 3988 => b"1111111010111",  3989 => b"1111111010111",  3990 => b"1111111010111",  3991 => b"1111111011000",
 3992 => b"1111111011000",  3993 => b"1111111011001",  3994 => b"1111111011001",  3995 => b"1111111011001",
 3996 => b"1111111011010",  3997 => b"1111111011010",  3998 => b"1111111011010",  3999 => b"1111111011011",
 4000 => b"1111111011011",  4001 => b"1111111011100",  4002 => b"1111111011100",  4003 => b"1111111011100",
 4004 => b"1111111011101",  4005 => b"1111111011101",  4006 => b"1111111011110",  4007 => b"1111111011110",
 4008 => b"1111111011110",  4009 => b"1111111011111",  4010 => b"1111111011111",  4011 => b"1111111011111",
 4012 => b"1111111100000",  4013 => b"1111111100000",  4014 => b"1111111100001",  4015 => b"1111111100001",
 4016 => b"1111111100001",  4017 => b"1111111100010",  4018 => b"1111111100010",  4019 => b"1111111100011",
 4020 => b"1111111100011",  4021 => b"1111111100011",  4022 => b"1111111100100",  4023 => b"1111111100100",
 4024 => b"1111111100101",  4025 => b"1111111100101",  4026 => b"1111111100101",  4027 => b"1111111100110",
 4028 => b"1111111100110",  4029 => b"1111111100110",  4030 => b"1111111100111",  4031 => b"1111111100111",
 4032 => b"1111111101000",  4033 => b"1111111101000",  4034 => b"1111111101000",  4035 => b"1111111101001",
 4036 => b"1111111101001",  4037 => b"1111111101010",  4038 => b"1111111101010",  4039 => b"1111111101010",
 4040 => b"1111111101011",  4041 => b"1111111101011",  4042 => b"1111111101100",  4043 => b"1111111101100",
 4044 => b"1111111101100",  4045 => b"1111111101101",  4046 => b"1111111101101",  4047 => b"1111111101101",
 4048 => b"1111111101110",  4049 => b"1111111101110",  4050 => b"1111111101111",  4051 => b"1111111101111",
 4052 => b"1111111101111",  4053 => b"1111111110000",  4054 => b"1111111110000",  4055 => b"1111111110001",
 4056 => b"1111111110001",  4057 => b"1111111110001",  4058 => b"1111111110010",  4059 => b"1111111110010",
 4060 => b"1111111110011",  4061 => b"1111111110011",  4062 => b"1111111110011",  4063 => b"1111111110100",
 4064 => b"1111111110100",  4065 => b"1111111110101",  4066 => b"1111111110101",  4067 => b"1111111110101",
 4068 => b"1111111110110",  4069 => b"1111111110110",  4070 => b"1111111110110",  4071 => b"1111111110111",
 4072 => b"1111111110111",  4073 => b"1111111111000",  4074 => b"1111111111000",  4075 => b"1111111111000",
 4076 => b"1111111111001",  4077 => b"1111111111001",  4078 => b"1111111111010",  4079 => b"1111111111010",
 4080 => b"1111111111010",  4081 => b"1111111111011",  4082 => b"1111111111011",  4083 => b"1111111111100",
 4084 => b"1111111111100",  4085 => b"1111111111100",  4086 => b"1111111111101",  4087 => b"1111111111101",
 4088 => b"1111111111110",  4089 => b"1111111111110",  4090 => b"1111111111110",  4091 => b"1111111111111",
 4092 => b"1111111111111",  4093 => b"0000000000000",  4094 => b"0000000000000",  4095 => b"0000000000000",
 4096 => b"0000000000000",  4097 => b"0000000000000",  4098 => b"0000000000000",  4099 => b"0000000000001",
 4100 => b"0000000000001",  4101 => b"0000000000010",  4102 => b"0000000000010",  4103 => b"0000000000010",
 4104 => b"0000000000011",  4105 => b"0000000000011",  4106 => b"0000000000100",  4107 => b"0000000000100",
 4108 => b"0000000000100",  4109 => b"0000000000101",  4110 => b"0000000000101",  4111 => b"0000000000110",
 4112 => b"0000000000110",  4113 => b"0000000000110",  4114 => b"0000000000111",  4115 => b"0000000000111",
 4116 => b"0000000001000",  4117 => b"0000000001000",  4118 => b"0000000001000",  4119 => b"0000000001001",
 4120 => b"0000000001001",  4121 => b"0000000001010",  4122 => b"0000000001010",  4123 => b"0000000001010",
 4124 => b"0000000001011",  4125 => b"0000000001011",  4126 => b"0000000001011",  4127 => b"0000000001100",
 4128 => b"0000000001100",  4129 => b"0000000001101",  4130 => b"0000000001101",  4131 => b"0000000001101",
 4132 => b"0000000001110",  4133 => b"0000000001110",  4134 => b"0000000001111",  4135 => b"0000000001111",
 4136 => b"0000000001111",  4137 => b"0000000010000",  4138 => b"0000000010000",  4139 => b"0000000010001",
 4140 => b"0000000010001",  4141 => b"0000000010001",  4142 => b"0000000010010",  4143 => b"0000000010010",
 4144 => b"0000000010011",  4145 => b"0000000010011",  4146 => b"0000000010011",  4147 => b"0000000010100",
 4148 => b"0000000010100",  4149 => b"0000000010100",  4150 => b"0000000010101",  4151 => b"0000000010101",
 4152 => b"0000000010110",  4153 => b"0000000010110",  4154 => b"0000000010110",  4155 => b"0000000010111",
 4156 => b"0000000010111",  4157 => b"0000000011000",  4158 => b"0000000011000",  4159 => b"0000000011000",
 4160 => b"0000000011001",  4161 => b"0000000011001",  4162 => b"0000000011010",  4163 => b"0000000011010",
 4164 => b"0000000011010",  4165 => b"0000000011011",  4166 => b"0000000011011",  4167 => b"0000000011011",
 4168 => b"0000000011100",  4169 => b"0000000011100",  4170 => b"0000000011101",  4171 => b"0000000011101",
 4172 => b"0000000011101",  4173 => b"0000000011110",  4174 => b"0000000011110",  4175 => b"0000000011111",
 4176 => b"0000000011111",  4177 => b"0000000011111",  4178 => b"0000000100000",  4179 => b"0000000100000",
 4180 => b"0000000100001",  4181 => b"0000000100001",  4182 => b"0000000100001",  4183 => b"0000000100010",
 4184 => b"0000000100010",  4185 => b"0000000100010",  4186 => b"0000000100011",  4187 => b"0000000100011",
 4188 => b"0000000100100",  4189 => b"0000000100100",  4190 => b"0000000100100",  4191 => b"0000000100101",
 4192 => b"0000000100101",  4193 => b"0000000100110",  4194 => b"0000000100110",  4195 => b"0000000100110",
 4196 => b"0000000100111",  4197 => b"0000000100111",  4198 => b"0000000100111",  4199 => b"0000000101000",
 4200 => b"0000000101000",  4201 => b"0000000101001",  4202 => b"0000000101001",  4203 => b"0000000101001",
 4204 => b"0000000101010",  4205 => b"0000000101010",  4206 => b"0000000101011",  4207 => b"0000000101011",
 4208 => b"0000000101011",  4209 => b"0000000101100",  4210 => b"0000000101100",  4211 => b"0000000101100",
 4212 => b"0000000101101",  4213 => b"0000000101101",  4214 => b"0000000101110",  4215 => b"0000000101110",
 4216 => b"0000000101110",  4217 => b"0000000101111",  4218 => b"0000000101111",  4219 => b"0000000101111",
 4220 => b"0000000110000",  4221 => b"0000000110000",  4222 => b"0000000110001",  4223 => b"0000000110001",
 4224 => b"0000000110001",  4225 => b"0000000110010",  4226 => b"0000000110010",  4227 => b"0000000110011",
 4228 => b"0000000110011",  4229 => b"0000000110011",  4230 => b"0000000110100",  4231 => b"0000000110100",
 4232 => b"0000000110100",  4233 => b"0000000110101",  4234 => b"0000000110101",  4235 => b"0000000110110",
 4236 => b"0000000110110",  4237 => b"0000000110110",  4238 => b"0000000110111",  4239 => b"0000000110111",
 4240 => b"0000000110111",  4241 => b"0000000111000",  4242 => b"0000000111000",  4243 => b"0000000111001",
 4244 => b"0000000111001",  4245 => b"0000000111001",  4246 => b"0000000111010",  4247 => b"0000000111010",
 4248 => b"0000000111010",  4249 => b"0000000111011",  4250 => b"0000000111011",  4251 => b"0000000111100",
 4252 => b"0000000111100",  4253 => b"0000000111100",  4254 => b"0000000111101",  4255 => b"0000000111101",
 4256 => b"0000000111101",  4257 => b"0000000111110",  4258 => b"0000000111110",  4259 => b"0000000111111",
 4260 => b"0000000111111",  4261 => b"0000000111111",  4262 => b"0000001000000",  4263 => b"0000001000000",
 4264 => b"0000001000000",  4265 => b"0000001000001",  4266 => b"0000001000001",  4267 => b"0000001000010",
 4268 => b"0000001000010",  4269 => b"0000001000010",  4270 => b"0000001000011",  4271 => b"0000001000011",
 4272 => b"0000001000011",  4273 => b"0000001000100",  4274 => b"0000001000100",  4275 => b"0000001000100",
 4276 => b"0000001000101",  4277 => b"0000001000101",  4278 => b"0000001000110",  4279 => b"0000001000110",
 4280 => b"0000001000110",  4281 => b"0000001000111",  4282 => b"0000001000111",  4283 => b"0000001000111",
 4284 => b"0000001001000",  4285 => b"0000001001000",  4286 => b"0000001001000",  4287 => b"0000001001001",
 4288 => b"0000001001001",  4289 => b"0000001001010",  4290 => b"0000001001010",  4291 => b"0000001001010",
 4292 => b"0000001001011",  4293 => b"0000001001011",  4294 => b"0000001001011",  4295 => b"0000001001100",
 4296 => b"0000001001100",  4297 => b"0000001001100",  4298 => b"0000001001101",  4299 => b"0000001001101",
 4300 => b"0000001001110",  4301 => b"0000001001110",  4302 => b"0000001001110",  4303 => b"0000001001111",
 4304 => b"0000001001111",  4305 => b"0000001001111",  4306 => b"0000001010000",  4307 => b"0000001010000",
 4308 => b"0000001010000",  4309 => b"0000001010001",  4310 => b"0000001010001",  4311 => b"0000001010001",
 4312 => b"0000001010010",  4313 => b"0000001010010",  4314 => b"0000001010011",  4315 => b"0000001010011",
 4316 => b"0000001010011",  4317 => b"0000001010100",  4318 => b"0000001010100",  4319 => b"0000001010100",
 4320 => b"0000001010101",  4321 => b"0000001010101",  4322 => b"0000001010101",  4323 => b"0000001010110",
 4324 => b"0000001010110",  4325 => b"0000001010110",  4326 => b"0000001010111",  4327 => b"0000001010111",
 4328 => b"0000001010111",  4329 => b"0000001011000",  4330 => b"0000001011000",  4331 => b"0000001011000",
 4332 => b"0000001011001",  4333 => b"0000001011001",  4334 => b"0000001011010",  4335 => b"0000001011010",
 4336 => b"0000001011010",  4337 => b"0000001011011",  4338 => b"0000001011011",  4339 => b"0000001011011",
 4340 => b"0000001011100",  4341 => b"0000001011100",  4342 => b"0000001011100",  4343 => b"0000001011101",
 4344 => b"0000001011101",  4345 => b"0000001011101",  4346 => b"0000001011110",  4347 => b"0000001011110",
 4348 => b"0000001011110",  4349 => b"0000001011111",  4350 => b"0000001011111",  4351 => b"0000001011111",
 4352 => b"0000001100000",  4353 => b"0000001100000",  4354 => b"0000001100000",  4355 => b"0000001100001",
 4356 => b"0000001100001",  4357 => b"0000001100001",  4358 => b"0000001100010",  4359 => b"0000001100010",
 4360 => b"0000001100010",  4361 => b"0000001100011",  4362 => b"0000001100011",  4363 => b"0000001100011",
 4364 => b"0000001100100",  4365 => b"0000001100100",  4366 => b"0000001100100",  4367 => b"0000001100101",
 4368 => b"0000001100101",  4369 => b"0000001100101",  4370 => b"0000001100110",  4371 => b"0000001100110",
 4372 => b"0000001100110",  4373 => b"0000001100111",  4374 => b"0000001100111",  4375 => b"0000001100111",
 4376 => b"0000001101000",  4377 => b"0000001101000",  4378 => b"0000001101000",  4379 => b"0000001101001",
 4380 => b"0000001101001",  4381 => b"0000001101001",  4382 => b"0000001101010",  4383 => b"0000001101010",
 4384 => b"0000001101010",  4385 => b"0000001101011",  4386 => b"0000001101011",  4387 => b"0000001101011",
 4388 => b"0000001101100",  4389 => b"0000001101100",  4390 => b"0000001101100",  4391 => b"0000001101101",
 4392 => b"0000001101101",  4393 => b"0000001101101",  4394 => b"0000001101110",  4395 => b"0000001101110",
 4396 => b"0000001101110",  4397 => b"0000001101111",  4398 => b"0000001101111",  4399 => b"0000001101111",
 4400 => b"0000001110000",  4401 => b"0000001110000",  4402 => b"0000001110000",  4403 => b"0000001110001",
 4404 => b"0000001110001",  4405 => b"0000001110001",  4406 => b"0000001110001",  4407 => b"0000001110010",
 4408 => b"0000001110010",  4409 => b"0000001110010",  4410 => b"0000001110011",  4411 => b"0000001110011",
 4412 => b"0000001110011",  4413 => b"0000001110100",  4414 => b"0000001110100",  4415 => b"0000001110100",
 4416 => b"0000001110101",  4417 => b"0000001110101",  4418 => b"0000001110101",  4419 => b"0000001110110",
 4420 => b"0000001110110",  4421 => b"0000001110110",  4422 => b"0000001110110",  4423 => b"0000001110111",
 4424 => b"0000001110111",  4425 => b"0000001110111",  4426 => b"0000001111000",  4427 => b"0000001111000",
 4428 => b"0000001111000",  4429 => b"0000001111001",  4430 => b"0000001111001",  4431 => b"0000001111001",
 4432 => b"0000001111010",  4433 => b"0000001111010",  4434 => b"0000001111010",  4435 => b"0000001111010",
 4436 => b"0000001111011",  4437 => b"0000001111011",  4438 => b"0000001111011",  4439 => b"0000001111100",
 4440 => b"0000001111100",  4441 => b"0000001111100",  4442 => b"0000001111101",  4443 => b"0000001111101",
 4444 => b"0000001111101",  4445 => b"0000001111101",  4446 => b"0000001111110",  4447 => b"0000001111110",
 4448 => b"0000001111110",  4449 => b"0000001111111",  4450 => b"0000001111111",  4451 => b"0000001111111",
 4452 => b"0000001111111",  4453 => b"0000010000000",  4454 => b"0000010000000",  4455 => b"0000010000000",
 4456 => b"0000010000001",  4457 => b"0000010000001",  4458 => b"0000010000001",  4459 => b"0000010000010",
 4460 => b"0000010000010",  4461 => b"0000010000010",  4462 => b"0000010000010",  4463 => b"0000010000011",
 4464 => b"0000010000011",  4465 => b"0000010000011",  4466 => b"0000010000100",  4467 => b"0000010000100",
 4468 => b"0000010000100",  4469 => b"0000010000100",  4470 => b"0000010000101",  4471 => b"0000010000101",
 4472 => b"0000010000101",  4473 => b"0000010000110",  4474 => b"0000010000110",  4475 => b"0000010000110",
 4476 => b"0000010000110",  4477 => b"0000010000111",  4478 => b"0000010000111",  4479 => b"0000010000111",
 4480 => b"0000010000111",  4481 => b"0000010001000",  4482 => b"0000010001000",  4483 => b"0000010001000",
 4484 => b"0000010001001",  4485 => b"0000010001001",  4486 => b"0000010001001",  4487 => b"0000010001001",
 4488 => b"0000010001010",  4489 => b"0000010001010",  4490 => b"0000010001010",  4491 => b"0000010001010",
 4492 => b"0000010001011",  4493 => b"0000010001011",  4494 => b"0000010001011",  4495 => b"0000010001100",
 4496 => b"0000010001100",  4497 => b"0000010001100",  4498 => b"0000010001100",  4499 => b"0000010001101",
 4500 => b"0000010001101",  4501 => b"0000010001101",  4502 => b"0000010001101",  4503 => b"0000010001110",
 4504 => b"0000010001110",  4505 => b"0000010001110",  4506 => b"0000010001110",  4507 => b"0000010001111",
 4508 => b"0000010001111",  4509 => b"0000010001111",  4510 => b"0000010010000",  4511 => b"0000010010000",
 4512 => b"0000010010000",  4513 => b"0000010010000",  4514 => b"0000010010001",  4515 => b"0000010010001",
 4516 => b"0000010010001",  4517 => b"0000010010001",  4518 => b"0000010010010",  4519 => b"0000010010010",
 4520 => b"0000010010010",  4521 => b"0000010010010",  4522 => b"0000010010011",  4523 => b"0000010010011",
 4524 => b"0000010010011",  4525 => b"0000010010011",  4526 => b"0000010010100",  4527 => b"0000010010100",
 4528 => b"0000010010100",  4529 => b"0000010010100",  4530 => b"0000010010101",  4531 => b"0000010010101",
 4532 => b"0000010010101",  4533 => b"0000010010101",  4534 => b"0000010010110",  4535 => b"0000010010110",
 4536 => b"0000010010110",  4537 => b"0000010010110",  4538 => b"0000010010111",  4539 => b"0000010010111",
 4540 => b"0000010010111",  4541 => b"0000010010111",  4542 => b"0000010010111",  4543 => b"0000010011000",
 4544 => b"0000010011000",  4545 => b"0000010011000",  4546 => b"0000010011000",  4547 => b"0000010011001",
 4548 => b"0000010011001",  4549 => b"0000010011001",  4550 => b"0000010011001",  4551 => b"0000010011010",
 4552 => b"0000010011010",  4553 => b"0000010011010",  4554 => b"0000010011010",  4555 => b"0000010011011",
 4556 => b"0000010011011",  4557 => b"0000010011011",  4558 => b"0000010011011",  4559 => b"0000010011011",
 4560 => b"0000010011100",  4561 => b"0000010011100",  4562 => b"0000010011100",  4563 => b"0000010011100",
 4564 => b"0000010011101",  4565 => b"0000010011101",  4566 => b"0000010011101",  4567 => b"0000010011101",
 4568 => b"0000010011101",  4569 => b"0000010011110",  4570 => b"0000010011110",  4571 => b"0000010011110",
 4572 => b"0000010011110",  4573 => b"0000010011111",  4574 => b"0000010011111",  4575 => b"0000010011111",
 4576 => b"0000010011111",  4577 => b"0000010011111",  4578 => b"0000010100000",  4579 => b"0000010100000",
 4580 => b"0000010100000",  4581 => b"0000010100000",  4582 => b"0000010100000",  4583 => b"0000010100001",
 4584 => b"0000010100001",  4585 => b"0000010100001",  4586 => b"0000010100001",  4587 => b"0000010100010",
 4588 => b"0000010100010",  4589 => b"0000010100010",  4590 => b"0000010100010",  4591 => b"0000010100010",
 4592 => b"0000010100011",  4593 => b"0000010100011",  4594 => b"0000010100011",  4595 => b"0000010100011",
 4596 => b"0000010100011",  4597 => b"0000010100100",  4598 => b"0000010100100",  4599 => b"0000010100100",
 4600 => b"0000010100100",  4601 => b"0000010100100",  4602 => b"0000010100101",  4603 => b"0000010100101",
 4604 => b"0000010100101",  4605 => b"0000010100101",  4606 => b"0000010100101",  4607 => b"0000010100110",
 4608 => b"0000010100110",  4609 => b"0000010100110",  4610 => b"0000010100110",  4611 => b"0000010100110",
 4612 => b"0000010100110",  4613 => b"0000010100111",  4614 => b"0000010100111",  4615 => b"0000010100111",
 4616 => b"0000010100111",  4617 => b"0000010100111",  4618 => b"0000010101000",  4619 => b"0000010101000",
 4620 => b"0000010101000",  4621 => b"0000010101000",  4622 => b"0000010101000",  4623 => b"0000010101001",
 4624 => b"0000010101001",  4625 => b"0000010101001",  4626 => b"0000010101001",  4627 => b"0000010101001",
 4628 => b"0000010101001",  4629 => b"0000010101010",  4630 => b"0000010101010",  4631 => b"0000010101010",
 4632 => b"0000010101010",  4633 => b"0000010101010",  4634 => b"0000010101010",  4635 => b"0000010101011",
 4636 => b"0000010101011",  4637 => b"0000010101011",  4638 => b"0000010101011",  4639 => b"0000010101011",
 4640 => b"0000010101011",  4641 => b"0000010101100",  4642 => b"0000010101100",  4643 => b"0000010101100",
 4644 => b"0000010101100",  4645 => b"0000010101100",  4646 => b"0000010101100",  4647 => b"0000010101101",
 4648 => b"0000010101101",  4649 => b"0000010101101",  4650 => b"0000010101101",  4651 => b"0000010101101",
 4652 => b"0000010101101",  4653 => b"0000010101110",  4654 => b"0000010101110",  4655 => b"0000010101110",
 4656 => b"0000010101110",  4657 => b"0000010101110",  4658 => b"0000010101110",  4659 => b"0000010101111",
 4660 => b"0000010101111",  4661 => b"0000010101111",  4662 => b"0000010101111",  4663 => b"0000010101111",
 4664 => b"0000010101111",  4665 => b"0000010101111",  4666 => b"0000010110000",  4667 => b"0000010110000",
 4668 => b"0000010110000",  4669 => b"0000010110000",  4670 => b"0000010110000",  4671 => b"0000010110000",
 4672 => b"0000010110000",  4673 => b"0000010110001",  4674 => b"0000010110001",  4675 => b"0000010110001",
 4676 => b"0000010110001",  4677 => b"0000010110001",  4678 => b"0000010110001",  4679 => b"0000010110001",
 4680 => b"0000010110010",  4681 => b"0000010110010",  4682 => b"0000010110010",  4683 => b"0000010110010",
 4684 => b"0000010110010",  4685 => b"0000010110010",  4686 => b"0000010110010",  4687 => b"0000010110011",
 4688 => b"0000010110011",  4689 => b"0000010110011",  4690 => b"0000010110011",  4691 => b"0000010110011",
 4692 => b"0000010110011",  4693 => b"0000010110011",  4694 => b"0000010110011",  4695 => b"0000010110100",
 4696 => b"0000010110100",  4697 => b"0000010110100",  4698 => b"0000010110100",  4699 => b"0000010110100",
 4700 => b"0000010110100",  4701 => b"0000010110100",  4702 => b"0000010110100",  4703 => b"0000010110100",
 4704 => b"0000010110101",  4705 => b"0000010110101",  4706 => b"0000010110101",  4707 => b"0000010110101",
 4708 => b"0000010110101",  4709 => b"0000010110101",  4710 => b"0000010110101",  4711 => b"0000010110101",
 4712 => b"0000010110110",  4713 => b"0000010110110",  4714 => b"0000010110110",  4715 => b"0000010110110",
 4716 => b"0000010110110",  4717 => b"0000010110110",  4718 => b"0000010110110",  4719 => b"0000010110110",
 4720 => b"0000010110110",  4721 => b"0000010110110",  4722 => b"0000010110111",  4723 => b"0000010110111",
 4724 => b"0000010110111",  4725 => b"0000010110111",  4726 => b"0000010110111",  4727 => b"0000010110111",
 4728 => b"0000010110111",  4729 => b"0000010110111",  4730 => b"0000010110111",  4731 => b"0000010110111",
 4732 => b"0000010111000",  4733 => b"0000010111000",  4734 => b"0000010111000",  4735 => b"0000010111000",
 4736 => b"0000010111000",  4737 => b"0000010111000",  4738 => b"0000010111000",  4739 => b"0000010111000",
 4740 => b"0000010111000",  4741 => b"0000010111000",  4742 => b"0000010111000",  4743 => b"0000010111001",
 4744 => b"0000010111001",  4745 => b"0000010111001",  4746 => b"0000010111001",  4747 => b"0000010111001",
 4748 => b"0000010111001",  4749 => b"0000010111001",  4750 => b"0000010111001",  4751 => b"0000010111001",
 4752 => b"0000010111001",  4753 => b"0000010111001",  4754 => b"0000010111001",  4755 => b"0000010111001",
 4756 => b"0000010111010",  4757 => b"0000010111010",  4758 => b"0000010111010",  4759 => b"0000010111010",
 4760 => b"0000010111010",  4761 => b"0000010111010",  4762 => b"0000010111010",  4763 => b"0000010111010",
 4764 => b"0000010111010",  4765 => b"0000010111010",  4766 => b"0000010111010",  4767 => b"0000010111010",
 4768 => b"0000010111010",  4769 => b"0000010111010",  4770 => b"0000010111010",  4771 => b"0000010111011",
 4772 => b"0000010111011",  4773 => b"0000010111011",  4774 => b"0000010111011",  4775 => b"0000010111011",
 4776 => b"0000010111011",  4777 => b"0000010111011",  4778 => b"0000010111011",  4779 => b"0000010111011",
 4780 => b"0000010111011",  4781 => b"0000010111011",  4782 => b"0000010111011",  4783 => b"0000010111011",
 4784 => b"0000010111011",  4785 => b"0000010111011",  4786 => b"0000010111011",  4787 => b"0000010111011",
 4788 => b"0000010111011",  4789 => b"0000010111011",  4790 => b"0000010111011",  4791 => b"0000010111100",
 4792 => b"0000010111100",  4793 => b"0000010111100",  4794 => b"0000010111100",  4795 => b"0000010111100",
 4796 => b"0000010111100",  4797 => b"0000010111100",  4798 => b"0000010111100",  4799 => b"0000010111100",
 4800 => b"0000010111100",  4801 => b"0000010111100",  4802 => b"0000010111100",  4803 => b"0000010111100",
 4804 => b"0000010111100",  4805 => b"0000010111100",  4806 => b"0000010111100",  4807 => b"0000010111100",
 4808 => b"0000010111100",  4809 => b"0000010111100",  4810 => b"0000010111100",  4811 => b"0000010111100",
 4812 => b"0000010111100",  4813 => b"0000010111100",  4814 => b"0000010111100",  4815 => b"0000010111100",
 4816 => b"0000010111100",  4817 => b"0000010111100",  4818 => b"0000010111100",  4819 => b"0000010111100",
 4820 => b"0000010111100",  4821 => b"0000010111100",  4822 => b"0000010111100",  4823 => b"0000010111100",
 4824 => b"0000010111100",  4825 => b"0000010111100",  4826 => b"0000010111100",  4827 => b"0000010111100",
 4828 => b"0000010111100",  4829 => b"0000010111100",  4830 => b"0000010111100",  4831 => b"0000010111100",
 4832 => b"0000010111100",  4833 => b"0000010111100",  4834 => b"0000010111100",  4835 => b"0000010111100",
 4836 => b"0000010111100",  4837 => b"0000010111100",  4838 => b"0000010111100",  4839 => b"0000010111100",
 4840 => b"0000010111100",  4841 => b"0000010111100",  4842 => b"0000010111100",  4843 => b"0000010111100",
 4844 => b"0000010111100",  4845 => b"0000010111100",  4846 => b"0000010111100",  4847 => b"0000010111100",
 4848 => b"0000010111100",  4849 => b"0000010111100",  4850 => b"0000010111100",  4851 => b"0000010111100",
 4852 => b"0000010111100",  4853 => b"0000010111100",  4854 => b"0000010111100",  4855 => b"0000010111100",
 4856 => b"0000010111100",  4857 => b"0000010111100",  4858 => b"0000010111100",  4859 => b"0000010111100",
 4860 => b"0000010111100",  4861 => b"0000010111100",  4862 => b"0000010111100",  4863 => b"0000010111100",
 4864 => b"0000010111100",  4865 => b"0000010111100",  4866 => b"0000010111100",  4867 => b"0000010111100",
 4868 => b"0000010111100",  4869 => b"0000010111100",  4870 => b"0000010111100",  4871 => b"0000010111100",
 4872 => b"0000010111100",  4873 => b"0000010111100",  4874 => b"0000010111100",  4875 => b"0000010111100",
 4876 => b"0000010111100",  4877 => b"0000010111100",  4878 => b"0000010111100",  4879 => b"0000010111100",
 4880 => b"0000010111100",  4881 => b"0000010111011",  4882 => b"0000010111011",  4883 => b"0000010111011",
 4884 => b"0000010111011",  4885 => b"0000010111011",  4886 => b"0000010111011",  4887 => b"0000010111011",
 4888 => b"0000010111011",  4889 => b"0000010111011",  4890 => b"0000010111011",  4891 => b"0000010111011",
 4892 => b"0000010111011",  4893 => b"0000010111011",  4894 => b"0000010111011",  4895 => b"0000010111011",
 4896 => b"0000010111011",  4897 => b"0000010111011",  4898 => b"0000010111011",  4899 => b"0000010111011",
 4900 => b"0000010111010",  4901 => b"0000010111010",  4902 => b"0000010111010",  4903 => b"0000010111010",
 4904 => b"0000010111010",  4905 => b"0000010111010",  4906 => b"0000010111010",  4907 => b"0000010111010",
 4908 => b"0000010111010",  4909 => b"0000010111010",  4910 => b"0000010111010",  4911 => b"0000010111010",
 4912 => b"0000010111010",  4913 => b"0000010111010",  4914 => b"0000010111010",  4915 => b"0000010111001",
 4916 => b"0000010111001",  4917 => b"0000010111001",  4918 => b"0000010111001",  4919 => b"0000010111001",
 4920 => b"0000010111001",  4921 => b"0000010111001",  4922 => b"0000010111001",  4923 => b"0000010111001",
 4924 => b"0000010111001",  4925 => b"0000010111001",  4926 => b"0000010111001",  4927 => b"0000010111000",
 4928 => b"0000010111000",  4929 => b"0000010111000",  4930 => b"0000010111000",  4931 => b"0000010111000",
 4932 => b"0000010111000",  4933 => b"0000010111000",  4934 => b"0000010111000",  4935 => b"0000010111000",
 4936 => b"0000010111000",  4937 => b"0000010111000",  4938 => b"0000010110111",  4939 => b"0000010110111",
 4940 => b"0000010110111",  4941 => b"0000010110111",  4942 => b"0000010110111",  4943 => b"0000010110111",
 4944 => b"0000010110111",  4945 => b"0000010110111",  4946 => b"0000010110111",  4947 => b"0000010110111",
 4948 => b"0000010110110",  4949 => b"0000010110110",  4950 => b"0000010110110",  4951 => b"0000010110110",
 4952 => b"0000010110110",  4953 => b"0000010110110",  4954 => b"0000010110110",  4955 => b"0000010110110",
 4956 => b"0000010110110",  4957 => b"0000010110101",  4958 => b"0000010110101",  4959 => b"0000010110101",
 4960 => b"0000010110101",  4961 => b"0000010110101",  4962 => b"0000010110101",  4963 => b"0000010110101",
 4964 => b"0000010110101",  4965 => b"0000010110100",  4966 => b"0000010110100",  4967 => b"0000010110100",
 4968 => b"0000010110100",  4969 => b"0000010110100",  4970 => b"0000010110100",  4971 => b"0000010110100",
 4972 => b"0000010110100",  4973 => b"0000010110011",  4974 => b"0000010110011",  4975 => b"0000010110011",
 4976 => b"0000010110011",  4977 => b"0000010110011",  4978 => b"0000010110011",  4979 => b"0000010110011",
 4980 => b"0000010110011",  4981 => b"0000010110010",  4982 => b"0000010110010",  4983 => b"0000010110010",
 4984 => b"0000010110010",  4985 => b"0000010110010",  4986 => b"0000010110010",  4987 => b"0000010110010",
 4988 => b"0000010110001",  4989 => b"0000010110001",  4990 => b"0000010110001",  4991 => b"0000010110001",
 4992 => b"0000010110001",  4993 => b"0000010110001",  4994 => b"0000010110000",  4995 => b"0000010110000",
 4996 => b"0000010110000",  4997 => b"0000010110000",  4998 => b"0000010110000",  4999 => b"0000010110000",
 5000 => b"0000010110000",  5001 => b"0000010101111",  5002 => b"0000010101111",  5003 => b"0000010101111",
 5004 => b"0000010101111",  5005 => b"0000010101111",  5006 => b"0000010101111",  5007 => b"0000010101110",
 5008 => b"0000010101110",  5009 => b"0000010101110",  5010 => b"0000010101110",  5011 => b"0000010101110",
 5012 => b"0000010101110",  5013 => b"0000010101101",  5014 => b"0000010101101",  5015 => b"0000010101101",
 5016 => b"0000010101101",  5017 => b"0000010101101",  5018 => b"0000010101101",  5019 => b"0000010101100",
 5020 => b"0000010101100",  5021 => b"0000010101100",  5022 => b"0000010101100",  5023 => b"0000010101100",
 5024 => b"0000010101011",  5025 => b"0000010101011",  5026 => b"0000010101011",  5027 => b"0000010101011",
 5028 => b"0000010101011",  5029 => b"0000010101010",  5030 => b"0000010101010",  5031 => b"0000010101010",
 5032 => b"0000010101010",  5033 => b"0000010101010",  5034 => b"0000010101010",  5035 => b"0000010101001",
 5036 => b"0000010101001",  5037 => b"0000010101001",  5038 => b"0000010101001",  5039 => b"0000010101001",
 5040 => b"0000010101000",  5041 => b"0000010101000",  5042 => b"0000010101000",  5043 => b"0000010101000",
 5044 => b"0000010101000",  5045 => b"0000010100111",  5046 => b"0000010100111",  5047 => b"0000010100111",
 5048 => b"0000010100111",  5049 => b"0000010100111",  5050 => b"0000010100110",  5051 => b"0000010100110",
 5052 => b"0000010100110",  5053 => b"0000010100110",  5054 => b"0000010100101",  5055 => b"0000010100101",
 5056 => b"0000010100101",  5057 => b"0000010100101",  5058 => b"0000010100101",  5059 => b"0000010100100",
 5060 => b"0000010100100",  5061 => b"0000010100100",  5062 => b"0000010100100",  5063 => b"0000010100100",
 5064 => b"0000010100011",  5065 => b"0000010100011",  5066 => b"0000010100011",  5067 => b"0000010100011",
 5068 => b"0000010100010",  5069 => b"0000010100010",  5070 => b"0000010100010",  5071 => b"0000010100010",
 5072 => b"0000010100010",  5073 => b"0000010100001",  5074 => b"0000010100001",  5075 => b"0000010100001",
 5076 => b"0000010100001",  5077 => b"0000010100000",  5078 => b"0000010100000",  5079 => b"0000010100000",
 5080 => b"0000010100000",  5081 => b"0000010011111",  5082 => b"0000010011111",  5083 => b"0000010011111",
 5084 => b"0000010011111",  5085 => b"0000010011110",  5086 => b"0000010011110",  5087 => b"0000010011110",
 5088 => b"0000010011110",  5089 => b"0000010011101",  5090 => b"0000010011101",  5091 => b"0000010011101",
 5092 => b"0000010011101",  5093 => b"0000010011100",  5094 => b"0000010011100",  5095 => b"0000010011100",
 5096 => b"0000010011100",  5097 => b"0000010011011",  5098 => b"0000010011011",  5099 => b"0000010011011",
 5100 => b"0000010011011",  5101 => b"0000010011010",  5102 => b"0000010011010",  5103 => b"0000010011010",
 5104 => b"0000010011010",  5105 => b"0000010011001",  5106 => b"0000010011001",  5107 => b"0000010011001",
 5108 => b"0000010011001",  5109 => b"0000010011000",  5110 => b"0000010011000",  5111 => b"0000010011000",
 5112 => b"0000010010111",  5113 => b"0000010010111",  5114 => b"0000010010111",  5115 => b"0000010010111",
 5116 => b"0000010010110",  5117 => b"0000010010110",  5118 => b"0000010010110",  5119 => b"0000010010110",
 5120 => b"0000010010101",  5121 => b"0000010010101",  5122 => b"0000010010101",  5123 => b"0000010010100",
 5124 => b"0000010010100",  5125 => b"0000010010100",  5126 => b"0000010010100",  5127 => b"0000010010011",
 5128 => b"0000010010011",  5129 => b"0000010010011",  5130 => b"0000010010010",  5131 => b"0000010010010",
 5132 => b"0000010010010",  5133 => b"0000010010010",  5134 => b"0000010010001",  5135 => b"0000010010001",
 5136 => b"0000010010001",  5137 => b"0000010010000",  5138 => b"0000010010000",  5139 => b"0000010010000",
 5140 => b"0000010010000",  5141 => b"0000010001111",  5142 => b"0000010001111",  5143 => b"0000010001111",
 5144 => b"0000010001110",  5145 => b"0000010001110",  5146 => b"0000010001110",  5147 => b"0000010001101",
 5148 => b"0000010001101",  5149 => b"0000010001101",  5150 => b"0000010001100",  5151 => b"0000010001100",
 5152 => b"0000010001100",  5153 => b"0000010001100",  5154 => b"0000010001011",  5155 => b"0000010001011",
 5156 => b"0000010001011",  5157 => b"0000010001010",  5158 => b"0000010001010",  5159 => b"0000010001010",
 5160 => b"0000010001001",  5161 => b"0000010001001",  5162 => b"0000010001001",  5163 => b"0000010001000",
 5164 => b"0000010001000",  5165 => b"0000010001000",  5166 => b"0000010000111",  5167 => b"0000010000111",
 5168 => b"0000010000111",  5169 => b"0000010000110",  5170 => b"0000010000110",  5171 => b"0000010000110",
 5172 => b"0000010000101",  5173 => b"0000010000101",  5174 => b"0000010000101",  5175 => b"0000010000100",
 5176 => b"0000010000100",  5177 => b"0000010000100",  5178 => b"0000010000011",  5179 => b"0000010000011",
 5180 => b"0000010000011",  5181 => b"0000010000010",  5182 => b"0000010000010",  5183 => b"0000010000010",
 5184 => b"0000010000001",  5185 => b"0000010000001",  5186 => b"0000010000001",  5187 => b"0000010000000",
 5188 => b"0000010000000",  5189 => b"0000010000000",  5190 => b"0000001111111",  5191 => b"0000001111111",
 5192 => b"0000001111111",  5193 => b"0000001111110",  5194 => b"0000001111110",  5195 => b"0000001111110",
 5196 => b"0000001111101",  5197 => b"0000001111101",  5198 => b"0000001111101",  5199 => b"0000001111100",
 5200 => b"0000001111100",  5201 => b"0000001111100",  5202 => b"0000001111011",  5203 => b"0000001111011",
 5204 => b"0000001111010",  5205 => b"0000001111010",  5206 => b"0000001111010",  5207 => b"0000001111001",
 5208 => b"0000001111001",  5209 => b"0000001111001",  5210 => b"0000001111000",  5211 => b"0000001111000",
 5212 => b"0000001111000",  5213 => b"0000001110111",  5214 => b"0000001110111",  5215 => b"0000001110110",
 5216 => b"0000001110110",  5217 => b"0000001110110",  5218 => b"0000001110101",  5219 => b"0000001110101",
 5220 => b"0000001110101",  5221 => b"0000001110100",  5222 => b"0000001110100",  5223 => b"0000001110011",
 5224 => b"0000001110011",  5225 => b"0000001110011",  5226 => b"0000001110010",  5227 => b"0000001110010",
 5228 => b"0000001110001",  5229 => b"0000001110001",  5230 => b"0000001110001",  5231 => b"0000001110000",
 5232 => b"0000001110000",  5233 => b"0000001110000",  5234 => b"0000001101111",  5235 => b"0000001101111",
 5236 => b"0000001101110",  5237 => b"0000001101110",  5238 => b"0000001101110",  5239 => b"0000001101101",
 5240 => b"0000001101101",  5241 => b"0000001101100",  5242 => b"0000001101100",  5243 => b"0000001101100",
 5244 => b"0000001101011",  5245 => b"0000001101011",  5246 => b"0000001101010",  5247 => b"0000001101010",
 5248 => b"0000001101010",  5249 => b"0000001101001",  5250 => b"0000001101001",  5251 => b"0000001101000",
 5252 => b"0000001101000",  5253 => b"0000001101000",  5254 => b"0000001100111",  5255 => b"0000001100111",
 5256 => b"0000001100110",  5257 => b"0000001100110",  5258 => b"0000001100110",  5259 => b"0000001100101",
 5260 => b"0000001100101",  5261 => b"0000001100100",  5262 => b"0000001100100",  5263 => b"0000001100011",
 5264 => b"0000001100011",  5265 => b"0000001100011",  5266 => b"0000001100010",  5267 => b"0000001100010",
 5268 => b"0000001100001",  5269 => b"0000001100001",  5270 => b"0000001100001",  5271 => b"0000001100000",
 5272 => b"0000001100000",  5273 => b"0000001011111",  5274 => b"0000001011111",  5275 => b"0000001011110",
 5276 => b"0000001011110",  5277 => b"0000001011110",  5278 => b"0000001011101",  5279 => b"0000001011101",
 5280 => b"0000001011100",  5281 => b"0000001011100",  5282 => b"0000001011011",  5283 => b"0000001011011",
 5284 => b"0000001011011",  5285 => b"0000001011010",  5286 => b"0000001011010",  5287 => b"0000001011001",
 5288 => b"0000001011001",  5289 => b"0000001011000",  5290 => b"0000001011000",  5291 => b"0000001010111",
 5292 => b"0000001010111",  5293 => b"0000001010111",  5294 => b"0000001010110",  5295 => b"0000001010110",
 5296 => b"0000001010101",  5297 => b"0000001010101",  5298 => b"0000001010100",  5299 => b"0000001010100",
 5300 => b"0000001010011",  5301 => b"0000001010011",  5302 => b"0000001010010",  5303 => b"0000001010010",
 5304 => b"0000001010010",  5305 => b"0000001010001",  5306 => b"0000001010001",  5307 => b"0000001010000",
 5308 => b"0000001010000",  5309 => b"0000001001111",  5310 => b"0000001001111",  5311 => b"0000001001110",
 5312 => b"0000001001110",  5313 => b"0000001001101",  5314 => b"0000001001101",  5315 => b"0000001001101",
 5316 => b"0000001001100",  5317 => b"0000001001100",  5318 => b"0000001001011",  5319 => b"0000001001011",
 5320 => b"0000001001010",  5321 => b"0000001001010",  5322 => b"0000001001001",  5323 => b"0000001001001",
 5324 => b"0000001001000",  5325 => b"0000001001000",  5326 => b"0000001000111",  5327 => b"0000001000111",
 5328 => b"0000001000110",  5329 => b"0000001000110",  5330 => b"0000001000101",  5331 => b"0000001000101",
 5332 => b"0000001000100",  5333 => b"0000001000100",  5334 => b"0000001000100",  5335 => b"0000001000011",
 5336 => b"0000001000011",  5337 => b"0000001000010",  5338 => b"0000001000010",  5339 => b"0000001000001",
 5340 => b"0000001000001",  5341 => b"0000001000000",  5342 => b"0000001000000",  5343 => b"0000000111111",
 5344 => b"0000000111111",  5345 => b"0000000111110",  5346 => b"0000000111110",  5347 => b"0000000111101",
 5348 => b"0000000111101",  5349 => b"0000000111100",  5350 => b"0000000111100",  5351 => b"0000000111011",
 5352 => b"0000000111011",  5353 => b"0000000111010",  5354 => b"0000000111010",  5355 => b"0000000111001",
 5356 => b"0000000111001",  5357 => b"0000000111000",  5358 => b"0000000111000",  5359 => b"0000000110111",
 5360 => b"0000000110111",  5361 => b"0000000110110",  5362 => b"0000000110110",  5363 => b"0000000110101",
 5364 => b"0000000110101",  5365 => b"0000000110100",  5366 => b"0000000110100",  5367 => b"0000000110011",
 5368 => b"0000000110011",  5369 => b"0000000110010",  5370 => b"0000000110010",  5371 => b"0000000110001",
 5372 => b"0000000110001",  5373 => b"0000000110000",  5374 => b"0000000110000",  5375 => b"0000000101111",
 5376 => b"0000000101110",  5377 => b"0000000101110",  5378 => b"0000000101101",  5379 => b"0000000101101",
 5380 => b"0000000101100",  5381 => b"0000000101100",  5382 => b"0000000101011",  5383 => b"0000000101011",
 5384 => b"0000000101010",  5385 => b"0000000101010",  5386 => b"0000000101001",  5387 => b"0000000101001",
 5388 => b"0000000101000",  5389 => b"0000000101000",  5390 => b"0000000100111",  5391 => b"0000000100111",
 5392 => b"0000000100110",  5393 => b"0000000100110",  5394 => b"0000000100101",  5395 => b"0000000100100",
 5396 => b"0000000100100",  5397 => b"0000000100011",  5398 => b"0000000100011",  5399 => b"0000000100010",
 5400 => b"0000000100010",  5401 => b"0000000100001",  5402 => b"0000000100001",  5403 => b"0000000100000",
 5404 => b"0000000100000",  5405 => b"0000000011111",  5406 => b"0000000011111",  5407 => b"0000000011110",
 5408 => b"0000000011101",  5409 => b"0000000011101",  5410 => b"0000000011100",  5411 => b"0000000011100",
 5412 => b"0000000011011",  5413 => b"0000000011011",  5414 => b"0000000011010",  5415 => b"0000000011010",
 5416 => b"0000000011001",  5417 => b"0000000011000",  5418 => b"0000000011000",  5419 => b"0000000010111",
 5420 => b"0000000010111",  5421 => b"0000000010110",  5422 => b"0000000010110",  5423 => b"0000000010101",
 5424 => b"0000000010101",  5425 => b"0000000010100",  5426 => b"0000000010011",  5427 => b"0000000010011",
 5428 => b"0000000010010",  5429 => b"0000000010010",  5430 => b"0000000010001",  5431 => b"0000000010001",
 5432 => b"0000000010000",  5433 => b"0000000001111",  5434 => b"0000000001111",  5435 => b"0000000001110",
 5436 => b"0000000001110",  5437 => b"0000000001101",  5438 => b"0000000001101",  5439 => b"0000000001100",
 5440 => b"0000000001100",  5441 => b"0000000001011",  5442 => b"0000000001010",  5443 => b"0000000001010",
 5444 => b"0000000001001",  5445 => b"0000000001001",  5446 => b"0000000001000",  5447 => b"0000000000111",
 5448 => b"0000000000111",  5449 => b"0000000000110",  5450 => b"0000000000110",  5451 => b"0000000000101",
 5452 => b"0000000000101",  5453 => b"0000000000100",  5454 => b"0000000000011",  5455 => b"0000000000011",
 5456 => b"0000000000010",  5457 => b"0000000000010",  5458 => b"0000000000001",  5459 => b"0000000000000",
 5460 => b"0000000000000",  5461 => b"0000000000000",  5462 => b"0000000000000",  5463 => b"1111111111111",
 5464 => b"1111111111111",  5465 => b"1111111111110",  5466 => b"1111111111101",  5467 => b"1111111111101",
 5468 => b"1111111111100",  5469 => b"1111111111100",  5470 => b"1111111111011",  5471 => b"1111111111010",
 5472 => b"1111111111010",  5473 => b"1111111111001",  5474 => b"1111111111001",  5475 => b"1111111111000",
 5476 => b"1111111110111",  5477 => b"1111111110111",  5478 => b"1111111110110",  5479 => b"1111111110110",
 5480 => b"1111111110101",  5481 => b"1111111110100",  5482 => b"1111111110100",  5483 => b"1111111110011",
 5484 => b"1111111110011",  5485 => b"1111111110010",  5486 => b"1111111110001",  5487 => b"1111111110001",
 5488 => b"1111111110000",  5489 => b"1111111101111",  5490 => b"1111111101111",  5491 => b"1111111101110",
 5492 => b"1111111101110",  5493 => b"1111111101101",  5494 => b"1111111101100",  5495 => b"1111111101100",
 5496 => b"1111111101011",  5497 => b"1111111101011",  5498 => b"1111111101010",  5499 => b"1111111101001",
 5500 => b"1111111101001",  5501 => b"1111111101000",  5502 => b"1111111100111",  5503 => b"1111111100111",
 5504 => b"1111111100110",  5505 => b"1111111100110",  5506 => b"1111111100101",  5507 => b"1111111100100",
 5508 => b"1111111100100",  5509 => b"1111111100011",  5510 => b"1111111100011",  5511 => b"1111111100010",
 5512 => b"1111111100001",  5513 => b"1111111100001",  5514 => b"1111111100000",  5515 => b"1111111011111",
 5516 => b"1111111011111",  5517 => b"1111111011110",  5518 => b"1111111011101",  5519 => b"1111111011101",
 5520 => b"1111111011100",  5521 => b"1111111011100",  5522 => b"1111111011011",  5523 => b"1111111011010",
 5524 => b"1111111011010",  5525 => b"1111111011001",  5526 => b"1111111011000",  5527 => b"1111111011000",
 5528 => b"1111111010111",  5529 => b"1111111010110",  5530 => b"1111111010110",  5531 => b"1111111010101",
 5532 => b"1111111010101",  5533 => b"1111111010100",  5534 => b"1111111010011",  5535 => b"1111111010011",
 5536 => b"1111111010010",  5537 => b"1111111010001",  5538 => b"1111111010001",  5539 => b"1111111010000",
 5540 => b"1111111001111",  5541 => b"1111111001111",  5542 => b"1111111001110",  5543 => b"1111111001101",
 5544 => b"1111111001101",  5545 => b"1111111001100",  5546 => b"1111111001011",  5547 => b"1111111001011",
 5548 => b"1111111001010",  5549 => b"1111111001010",  5550 => b"1111111001001",  5551 => b"1111111001000",
 5552 => b"1111111001000",  5553 => b"1111111000111",  5554 => b"1111111000110",  5555 => b"1111111000110",
 5556 => b"1111111000101",  5557 => b"1111111000100",  5558 => b"1111111000100",  5559 => b"1111111000011",
 5560 => b"1111111000010",  5561 => b"1111111000010",  5562 => b"1111111000001",  5563 => b"1111111000000",
 5564 => b"1111111000000",  5565 => b"1111110111111",  5566 => b"1111110111110",  5567 => b"1111110111110",
 5568 => b"1111110111101",  5569 => b"1111110111100",  5570 => b"1111110111100",  5571 => b"1111110111011",
 5572 => b"1111110111010",  5573 => b"1111110111010",  5574 => b"1111110111001",  5575 => b"1111110111000",
 5576 => b"1111110111000",  5577 => b"1111110110111",  5578 => b"1111110110110",  5579 => b"1111110110110",
 5580 => b"1111110110101",  5581 => b"1111110110100",  5582 => b"1111110110100",  5583 => b"1111110110011",
 5584 => b"1111110110010",  5585 => b"1111110110010",  5586 => b"1111110110001",  5587 => b"1111110110000",
 5588 => b"1111110110000",  5589 => b"1111110101111",  5590 => b"1111110101110",  5591 => b"1111110101101",
 5592 => b"1111110101101",  5593 => b"1111110101100",  5594 => b"1111110101011",  5595 => b"1111110101011",
 5596 => b"1111110101010",  5597 => b"1111110101001",  5598 => b"1111110101001",  5599 => b"1111110101000",
 5600 => b"1111110100111",  5601 => b"1111110100111",  5602 => b"1111110100110",  5603 => b"1111110100101",
 5604 => b"1111110100101",  5605 => b"1111110100100",  5606 => b"1111110100011",  5607 => b"1111110100010",
 5608 => b"1111110100010",  5609 => b"1111110100001",  5610 => b"1111110100000",  5611 => b"1111110100000",
 5612 => b"1111110011111",  5613 => b"1111110011110",  5614 => b"1111110011110",  5615 => b"1111110011101",
 5616 => b"1111110011100",  5617 => b"1111110011100",  5618 => b"1111110011011",  5619 => b"1111110011010",
 5620 => b"1111110011001",  5621 => b"1111110011001",  5622 => b"1111110011000",  5623 => b"1111110010111",
 5624 => b"1111110010111",  5625 => b"1111110010110",  5626 => b"1111110010101",  5627 => b"1111110010101",
 5628 => b"1111110010100",  5629 => b"1111110010011",  5630 => b"1111110010010",  5631 => b"1111110010010",
 5632 => b"1111110010001",  5633 => b"1111110010000",  5634 => b"1111110010000",  5635 => b"1111110001111",
 5636 => b"1111110001110",  5637 => b"1111110001101",  5638 => b"1111110001101",  5639 => b"1111110001100",
 5640 => b"1111110001011",  5641 => b"1111110001011",  5642 => b"1111110001010",  5643 => b"1111110001001",
 5644 => b"1111110001001",  5645 => b"1111110001000",  5646 => b"1111110000111",  5647 => b"1111110000110",
 5648 => b"1111110000110",  5649 => b"1111110000101",  5650 => b"1111110000100",  5651 => b"1111110000100",
 5652 => b"1111110000011",  5653 => b"1111110000010",  5654 => b"1111110000001",  5655 => b"1111110000001",
 5656 => b"1111110000000",  5657 => b"1111101111111",  5658 => b"1111101111110",  5659 => b"1111101111110",
 5660 => b"1111101111101",  5661 => b"1111101111100",  5662 => b"1111101111100",  5663 => b"1111101111011",
 5664 => b"1111101111010",  5665 => b"1111101111001",  5666 => b"1111101111001",  5667 => b"1111101111000",
 5668 => b"1111101110111",  5669 => b"1111101110111",  5670 => b"1111101110110",  5671 => b"1111101110101",
 5672 => b"1111101110100",  5673 => b"1111101110100",  5674 => b"1111101110011",  5675 => b"1111101110010",
 5676 => b"1111101110001",  5677 => b"1111101110001",  5678 => b"1111101110000",  5679 => b"1111101101111",
 5680 => b"1111101101110",  5681 => b"1111101101110",  5682 => b"1111101101101",  5683 => b"1111101101100",
 5684 => b"1111101101100",  5685 => b"1111101101011",  5686 => b"1111101101010",  5687 => b"1111101101001",
 5688 => b"1111101101001",  5689 => b"1111101101000",  5690 => b"1111101100111",  5691 => b"1111101100110",
 5692 => b"1111101100110",  5693 => b"1111101100101",  5694 => b"1111101100100",  5695 => b"1111101100011",
 5696 => b"1111101100011",  5697 => b"1111101100010",  5698 => b"1111101100001",  5699 => b"1111101100001",
 5700 => b"1111101100000",  5701 => b"1111101011111",  5702 => b"1111101011110",  5703 => b"1111101011110",
 5704 => b"1111101011101",  5705 => b"1111101011100",  5706 => b"1111101011011",  5707 => b"1111101011011",
 5708 => b"1111101011010",  5709 => b"1111101011001",  5710 => b"1111101011000",  5711 => b"1111101011000",
 5712 => b"1111101010111",  5713 => b"1111101010110",  5714 => b"1111101010101",  5715 => b"1111101010101",
 5716 => b"1111101010100",  5717 => b"1111101010011",  5718 => b"1111101010010",  5719 => b"1111101010010",
 5720 => b"1111101010001",  5721 => b"1111101010000",  5722 => b"1111101001111",  5723 => b"1111101001111",
 5724 => b"1111101001110",  5725 => b"1111101001101",  5726 => b"1111101001100",  5727 => b"1111101001100",
 5728 => b"1111101001011",  5729 => b"1111101001010",  5730 => b"1111101001001",  5731 => b"1111101001001",
 5732 => b"1111101001000",  5733 => b"1111101000111",  5734 => b"1111101000110",  5735 => b"1111101000110",
 5736 => b"1111101000101",  5737 => b"1111101000100",  5738 => b"1111101000011",  5739 => b"1111101000010",
 5740 => b"1111101000010",  5741 => b"1111101000001",  5742 => b"1111101000000",  5743 => b"1111100111111",
 5744 => b"1111100111111",  5745 => b"1111100111110",  5746 => b"1111100111101",  5747 => b"1111100111100",
 5748 => b"1111100111100",  5749 => b"1111100111011",  5750 => b"1111100111010",  5751 => b"1111100111001",
 5752 => b"1111100111001",  5753 => b"1111100111000",  5754 => b"1111100110111",  5755 => b"1111100110110",
 5756 => b"1111100110110",  5757 => b"1111100110101",  5758 => b"1111100110100",  5759 => b"1111100110011",
 5760 => b"1111100110010",  5761 => b"1111100110010",  5762 => b"1111100110001",  5763 => b"1111100110000",
 5764 => b"1111100101111",  5765 => b"1111100101111",  5766 => b"1111100101110",  5767 => b"1111100101101",
 5768 => b"1111100101100",  5769 => b"1111100101100",  5770 => b"1111100101011",  5771 => b"1111100101010",
 5772 => b"1111100101001",  5773 => b"1111100101000",  5774 => b"1111100101000",  5775 => b"1111100100111",
 5776 => b"1111100100110",  5777 => b"1111100100101",  5778 => b"1111100100101",  5779 => b"1111100100100",
 5780 => b"1111100100011",  5781 => b"1111100100010",  5782 => b"1111100100001",  5783 => b"1111100100001",
 5784 => b"1111100100000",  5785 => b"1111100011111",  5786 => b"1111100011110",  5787 => b"1111100011110",
 5788 => b"1111100011101",  5789 => b"1111100011100",  5790 => b"1111100011011",  5791 => b"1111100011010",
 5792 => b"1111100011010",  5793 => b"1111100011001",  5794 => b"1111100011000",  5795 => b"1111100010111",
 5796 => b"1111100010111",  5797 => b"1111100010110",  5798 => b"1111100010101",  5799 => b"1111100010100",
 5800 => b"1111100010011",  5801 => b"1111100010011",  5802 => b"1111100010010",  5803 => b"1111100010001",
 5804 => b"1111100010000",  5805 => b"1111100010000",  5806 => b"1111100001111",  5807 => b"1111100001110",
 5808 => b"1111100001101",  5809 => b"1111100001100",  5810 => b"1111100001100",  5811 => b"1111100001011",
 5812 => b"1111100001010",  5813 => b"1111100001001",  5814 => b"1111100001001",  5815 => b"1111100001000",
 5816 => b"1111100000111",  5817 => b"1111100000110",  5818 => b"1111100000101",  5819 => b"1111100000101",
 5820 => b"1111100000100",  5821 => b"1111100000011",  5822 => b"1111100000010",  5823 => b"1111100000001",
 5824 => b"1111100000001",  5825 => b"1111100000000",  5826 => b"1111011111111",  5827 => b"1111011111110",
 5828 => b"1111011111101",  5829 => b"1111011111101",  5830 => b"1111011111100",  5831 => b"1111011111011",
 5832 => b"1111011111010",  5833 => b"1111011111010",  5834 => b"1111011111001",  5835 => b"1111011111000",
 5836 => b"1111011110111",  5837 => b"1111011110110",  5838 => b"1111011110110",  5839 => b"1111011110101",
 5840 => b"1111011110100",  5841 => b"1111011110011",  5842 => b"1111011110010",  5843 => b"1111011110010",
 5844 => b"1111011110001",  5845 => b"1111011110000",  5846 => b"1111011101111",  5847 => b"1111011101110",
 5848 => b"1111011101110",  5849 => b"1111011101101",  5850 => b"1111011101100",  5851 => b"1111011101011",
 5852 => b"1111011101010",  5853 => b"1111011101010",  5854 => b"1111011101001",  5855 => b"1111011101000",
 5856 => b"1111011100111",  5857 => b"1111011100110",  5858 => b"1111011100110",  5859 => b"1111011100101",
 5860 => b"1111011100100",  5861 => b"1111011100011",  5862 => b"1111011100010",  5863 => b"1111011100010",
 5864 => b"1111011100001",  5865 => b"1111011100000",  5866 => b"1111011011111",  5867 => b"1111011011111",
 5868 => b"1111011011110",  5869 => b"1111011011101",  5870 => b"1111011011100",  5871 => b"1111011011011",
 5872 => b"1111011011011",  5873 => b"1111011011010",  5874 => b"1111011011001",  5875 => b"1111011011000",
 5876 => b"1111011010111",  5877 => b"1111011010111",  5878 => b"1111011010110",  5879 => b"1111011010101",
 5880 => b"1111011010100",  5881 => b"1111011010011",  5882 => b"1111011010011",  5883 => b"1111011010010",
 5884 => b"1111011010001",  5885 => b"1111011010000",  5886 => b"1111011001111",  5887 => b"1111011001110",
 5888 => b"1111011001110",  5889 => b"1111011001101",  5890 => b"1111011001100",  5891 => b"1111011001011",
 5892 => b"1111011001010",  5893 => b"1111011001010",  5894 => b"1111011001001",  5895 => b"1111011001000",
 5896 => b"1111011000111",  5897 => b"1111011000110",  5898 => b"1111011000110",  5899 => b"1111011000101",
 5900 => b"1111011000100",  5901 => b"1111011000011",  5902 => b"1111011000010",  5903 => b"1111011000010",
 5904 => b"1111011000001",  5905 => b"1111011000000",  5906 => b"1111010111111",  5907 => b"1111010111110",
 5908 => b"1111010111110",  5909 => b"1111010111101",  5910 => b"1111010111100",  5911 => b"1111010111011",
 5912 => b"1111010111010",  5913 => b"1111010111010",  5914 => b"1111010111001",  5915 => b"1111010111000",
 5916 => b"1111010110111",  5917 => b"1111010110110",  5918 => b"1111010110110",  5919 => b"1111010110101",
 5920 => b"1111010110100",  5921 => b"1111010110011",  5922 => b"1111010110010",  5923 => b"1111010110010",
 5924 => b"1111010110001",  5925 => b"1111010110000",  5926 => b"1111010101111",  5927 => b"1111010101110",
 5928 => b"1111010101101",  5929 => b"1111010101101",  5930 => b"1111010101100",  5931 => b"1111010101011",
 5932 => b"1111010101010",  5933 => b"1111010101001",  5934 => b"1111010101001",  5935 => b"1111010101000",
 5936 => b"1111010100111",  5937 => b"1111010100110",  5938 => b"1111010100101",  5939 => b"1111010100101",
 5940 => b"1111010100100",  5941 => b"1111010100011",  5942 => b"1111010100010",  5943 => b"1111010100001",
 5944 => b"1111010100001",  5945 => b"1111010100000",  5946 => b"1111010011111",  5947 => b"1111010011110",
 5948 => b"1111010011101",  5949 => b"1111010011101",  5950 => b"1111010011100",  5951 => b"1111010011011",
 5952 => b"1111010011010",  5953 => b"1111010011001",  5954 => b"1111010011000",  5955 => b"1111010011000",
 5956 => b"1111010010111",  5957 => b"1111010010110",  5958 => b"1111010010101",  5959 => b"1111010010100",
 5960 => b"1111010010100",  5961 => b"1111010010011",  5962 => b"1111010010010",  5963 => b"1111010010001",
 5964 => b"1111010010000",  5965 => b"1111010010000",  5966 => b"1111010001111",  5967 => b"1111010001110",
 5968 => b"1111010001101",  5969 => b"1111010001100",  5970 => b"1111010001100",  5971 => b"1111010001011",
 5972 => b"1111010001010",  5973 => b"1111010001001",  5974 => b"1111010001000",  5975 => b"1111010000111",
 5976 => b"1111010000111",  5977 => b"1111010000110",  5978 => b"1111010000101",  5979 => b"1111010000100",
 5980 => b"1111010000011",  5981 => b"1111010000011",  5982 => b"1111010000010",  5983 => b"1111010000001",
 5984 => b"1111010000000",  5985 => b"1111001111111",  5986 => b"1111001111111",  5987 => b"1111001111110",
 5988 => b"1111001111101",  5989 => b"1111001111100",  5990 => b"1111001111011",  5991 => b"1111001111010",
 5992 => b"1111001111010",  5993 => b"1111001111001",  5994 => b"1111001111000",  5995 => b"1111001110111",
 5996 => b"1111001110110",  5997 => b"1111001110110",  5998 => b"1111001110101",  5999 => b"1111001110100",
 6000 => b"1111001110011",  6001 => b"1111001110010",  6002 => b"1111001110010",  6003 => b"1111001110001",
 6004 => b"1111001110000",  6005 => b"1111001101111",  6006 => b"1111001101110",  6007 => b"1111001101110",
 6008 => b"1111001101101",  6009 => b"1111001101100",  6010 => b"1111001101011",  6011 => b"1111001101010",
 6012 => b"1111001101001",  6013 => b"1111001101001",  6014 => b"1111001101000",  6015 => b"1111001100111",
 6016 => b"1111001100110",  6017 => b"1111001100101",  6018 => b"1111001100101",  6019 => b"1111001100100",
 6020 => b"1111001100011",  6021 => b"1111001100010",  6022 => b"1111001100001",  6023 => b"1111001100001",
 6024 => b"1111001100000",  6025 => b"1111001011111",  6026 => b"1111001011110",  6027 => b"1111001011101",
 6028 => b"1111001011101",  6029 => b"1111001011100",  6030 => b"1111001011011",  6031 => b"1111001011010",
 6032 => b"1111001011001",  6033 => b"1111001011001",  6034 => b"1111001011000",  6035 => b"1111001010111",
 6036 => b"1111001010110",  6037 => b"1111001010101",  6038 => b"1111001010100",  6039 => b"1111001010100",
 6040 => b"1111001010011",  6041 => b"1111001010010",  6042 => b"1111001010001",  6043 => b"1111001010000",
 6044 => b"1111001010000",  6045 => b"1111001001111",  6046 => b"1111001001110",  6047 => b"1111001001101",
 6048 => b"1111001001100",  6049 => b"1111001001100",  6050 => b"1111001001011",  6051 => b"1111001001010",
 6052 => b"1111001001001",  6053 => b"1111001001000",  6054 => b"1111001001000",  6055 => b"1111001000111",
 6056 => b"1111001000110",  6057 => b"1111001000101",  6058 => b"1111001000100",  6059 => b"1111001000100",
 6060 => b"1111001000011",  6061 => b"1111001000010",  6062 => b"1111001000001",  6063 => b"1111001000000",
 6064 => b"1111001000000",  6065 => b"1111000111111",  6066 => b"1111000111110",  6067 => b"1111000111101",
 6068 => b"1111000111100",  6069 => b"1111000111100",  6070 => b"1111000111011",  6071 => b"1111000111010",
 6072 => b"1111000111001",  6073 => b"1111000111000",  6074 => b"1111000111000",  6075 => b"1111000110111",
 6076 => b"1111000110110",  6077 => b"1111000110101",  6078 => b"1111000110100",  6079 => b"1111000110100",
 6080 => b"1111000110011",  6081 => b"1111000110010",  6082 => b"1111000110001",  6083 => b"1111000110000",
 6084 => b"1111000110000",  6085 => b"1111000101111",  6086 => b"1111000101110",  6087 => b"1111000101101",
 6088 => b"1111000101100",  6089 => b"1111000101100",  6090 => b"1111000101011",  6091 => b"1111000101010",
 6092 => b"1111000101001",  6093 => b"1111000101000",  6094 => b"1111000101000",  6095 => b"1111000100111",
 6096 => b"1111000100110",  6097 => b"1111000100101",  6098 => b"1111000100100",  6099 => b"1111000100100",
 6100 => b"1111000100011",  6101 => b"1111000100010",  6102 => b"1111000100001",  6103 => b"1111000100000",
 6104 => b"1111000100000",  6105 => b"1111000011111",  6106 => b"1111000011110",  6107 => b"1111000011101",
 6108 => b"1111000011100",  6109 => b"1111000011100",  6110 => b"1111000011011",  6111 => b"1111000011010",
 6112 => b"1111000011001",  6113 => b"1111000011000",  6114 => b"1111000011000",  6115 => b"1111000010111",
 6116 => b"1111000010110",  6117 => b"1111000010101",  6118 => b"1111000010100",  6119 => b"1111000010100",
 6120 => b"1111000010011",  6121 => b"1111000010010",  6122 => b"1111000010001",  6123 => b"1111000010000",
 6124 => b"1111000010000",  6125 => b"1111000001111",  6126 => b"1111000001110",  6127 => b"1111000001101",
 6128 => b"1111000001101",  6129 => b"1111000001100",  6130 => b"1111000001011",  6131 => b"1111000001010",
 6132 => b"1111000001001",  6133 => b"1111000001001",  6134 => b"1111000001000",  6135 => b"1111000000111",
 6136 => b"1111000000110",  6137 => b"1111000000101",  6138 => b"1111000000101",  6139 => b"1111000000100",
 6140 => b"1111000000011",  6141 => b"1111000000010",  6142 => b"1111000000001",  6143 => b"1111000000001",
 6144 => b"1111000000000",  6145 => b"1110111111111",  6146 => b"1110111111110",  6147 => b"1110111111110",
 6148 => b"1110111111101",  6149 => b"1110111111100",  6150 => b"1110111111011",  6151 => b"1110111111010",
 6152 => b"1110111111010",  6153 => b"1110111111001",  6154 => b"1110111111000",  6155 => b"1110111110111",
 6156 => b"1110111110111",  6157 => b"1110111110110",  6158 => b"1110111110101",  6159 => b"1110111110100",
 6160 => b"1110111110011",  6161 => b"1110111110011",  6162 => b"1110111110010",  6163 => b"1110111110001",
 6164 => b"1110111110000",  6165 => b"1110111101111",  6166 => b"1110111101111",  6167 => b"1110111101110",
 6168 => b"1110111101101",  6169 => b"1110111101100",  6170 => b"1110111101100",  6171 => b"1110111101011",
 6172 => b"1110111101010",  6173 => b"1110111101001",  6174 => b"1110111101000",  6175 => b"1110111101000",
 6176 => b"1110111100111",  6177 => b"1110111100110",  6178 => b"1110111100101",  6179 => b"1110111100101",
 6180 => b"1110111100100",  6181 => b"1110111100011",  6182 => b"1110111100010",  6183 => b"1110111100010",
 6184 => b"1110111100001",  6185 => b"1110111100000",  6186 => b"1110111011111",  6187 => b"1110111011110",
 6188 => b"1110111011110",  6189 => b"1110111011101",  6190 => b"1110111011100",  6191 => b"1110111011011",
 6192 => b"1110111011011",  6193 => b"1110111011010",  6194 => b"1110111011001",  6195 => b"1110111011000",
 6196 => b"1110111011000",  6197 => b"1110111010111",  6198 => b"1110111010110",  6199 => b"1110111010101",
 6200 => b"1110111010100",  6201 => b"1110111010100",  6202 => b"1110111010011",  6203 => b"1110111010010",
 6204 => b"1110111010001",  6205 => b"1110111010001",  6206 => b"1110111010000",  6207 => b"1110111001111",
 6208 => b"1110111001110",  6209 => b"1110111001110",  6210 => b"1110111001101",  6211 => b"1110111001100",
 6212 => b"1110111001011",  6213 => b"1110111001011",  6214 => b"1110111001010",  6215 => b"1110111001001",
 6216 => b"1110111001000",  6217 => b"1110111001000",  6218 => b"1110111000111",  6219 => b"1110111000110",
 6220 => b"1110111000101",  6221 => b"1110111000100",  6222 => b"1110111000100",  6223 => b"1110111000011",
 6224 => b"1110111000010",  6225 => b"1110111000001",  6226 => b"1110111000001",  6227 => b"1110111000000",
 6228 => b"1110110111111",  6229 => b"1110110111110",  6230 => b"1110110111110",  6231 => b"1110110111101",
 6232 => b"1110110111100",  6233 => b"1110110111011",  6234 => b"1110110111011",  6235 => b"1110110111010",
 6236 => b"1110110111001",  6237 => b"1110110111000",  6238 => b"1110110111000",  6239 => b"1110110110111",
 6240 => b"1110110110110",  6241 => b"1110110110101",  6242 => b"1110110110101",  6243 => b"1110110110100",
 6244 => b"1110110110011",  6245 => b"1110110110010",  6246 => b"1110110110010",  6247 => b"1110110110001",
 6248 => b"1110110110000",  6249 => b"1110110101111",  6250 => b"1110110101111",  6251 => b"1110110101110",
 6252 => b"1110110101101",  6253 => b"1110110101101",  6254 => b"1110110101100",  6255 => b"1110110101011",
 6256 => b"1110110101010",  6257 => b"1110110101010",  6258 => b"1110110101001",  6259 => b"1110110101000",
 6260 => b"1110110100111",  6261 => b"1110110100111",  6262 => b"1110110100110",  6263 => b"1110110100101",
 6264 => b"1110110100100",  6265 => b"1110110100100",  6266 => b"1110110100011",  6267 => b"1110110100010",
 6268 => b"1110110100001",  6269 => b"1110110100001",  6270 => b"1110110100000",  6271 => b"1110110011111",
 6272 => b"1110110011111",  6273 => b"1110110011110",  6274 => b"1110110011101",  6275 => b"1110110011100",
 6276 => b"1110110011100",  6277 => b"1110110011011",  6278 => b"1110110011010",  6279 => b"1110110011001",
 6280 => b"1110110011001",  6281 => b"1110110011000",  6282 => b"1110110010111",  6283 => b"1110110010111",
 6284 => b"1110110010110",  6285 => b"1110110010101",  6286 => b"1110110010100",  6287 => b"1110110010100",
 6288 => b"1110110010011",  6289 => b"1110110010010",  6290 => b"1110110010001",  6291 => b"1110110010001",
 6292 => b"1110110010000",  6293 => b"1110110001111",  6294 => b"1110110001111",  6295 => b"1110110001110",
 6296 => b"1110110001101",  6297 => b"1110110001100",  6298 => b"1110110001100",  6299 => b"1110110001011",
 6300 => b"1110110001010",  6301 => b"1110110001010",  6302 => b"1110110001001",  6303 => b"1110110001000",
 6304 => b"1110110000111",  6305 => b"1110110000111",  6306 => b"1110110000110",  6307 => b"1110110000101",
 6308 => b"1110110000101",  6309 => b"1110110000100",  6310 => b"1110110000011",  6311 => b"1110110000010",
 6312 => b"1110110000010",  6313 => b"1110110000001",  6314 => b"1110110000000",  6315 => b"1110110000000",
 6316 => b"1110101111111",  6317 => b"1110101111110",  6318 => b"1110101111101",  6319 => b"1110101111101",
 6320 => b"1110101111100",  6321 => b"1110101111011",  6322 => b"1110101111011",  6323 => b"1110101111010",
 6324 => b"1110101111001",  6325 => b"1110101111001",  6326 => b"1110101111000",  6327 => b"1110101110111",
 6328 => b"1110101110110",  6329 => b"1110101110110",  6330 => b"1110101110101",  6331 => b"1110101110100",
 6332 => b"1110101110100",  6333 => b"1110101110011",  6334 => b"1110101110010",  6335 => b"1110101110010",
 6336 => b"1110101110001",  6337 => b"1110101110000",  6338 => b"1110101101111",  6339 => b"1110101101111",
 6340 => b"1110101101110",  6341 => b"1110101101101",  6342 => b"1110101101101",  6343 => b"1110101101100",
 6344 => b"1110101101011",  6345 => b"1110101101011",  6346 => b"1110101101010",  6347 => b"1110101101001",
 6348 => b"1110101101001",  6349 => b"1110101101000",  6350 => b"1110101100111",  6351 => b"1110101100111",
 6352 => b"1110101100110",  6353 => b"1110101100101",  6354 => b"1110101100101",  6355 => b"1110101100100",
 6356 => b"1110101100011",  6357 => b"1110101100010",  6358 => b"1110101100010",  6359 => b"1110101100001",
 6360 => b"1110101100000",  6361 => b"1110101100000",  6362 => b"1110101011111",  6363 => b"1110101011110",
 6364 => b"1110101011110",  6365 => b"1110101011101",  6366 => b"1110101011100",  6367 => b"1110101011100",
 6368 => b"1110101011011",  6369 => b"1110101011010",  6370 => b"1110101011010",  6371 => b"1110101011001",
 6372 => b"1110101011000",  6373 => b"1110101011000",  6374 => b"1110101010111",  6375 => b"1110101010110",
 6376 => b"1110101010110",  6377 => b"1110101010101",  6378 => b"1110101010100",  6379 => b"1110101010100",
 6380 => b"1110101010011",  6381 => b"1110101010010",  6382 => b"1110101010010",  6383 => b"1110101010001",
 6384 => b"1110101010000",  6385 => b"1110101010000",  6386 => b"1110101001111",  6387 => b"1110101001110",
 6388 => b"1110101001110",  6389 => b"1110101001101",  6390 => b"1110101001100",  6391 => b"1110101001100",
 6392 => b"1110101001011",  6393 => b"1110101001010",  6394 => b"1110101001010",  6395 => b"1110101001001",
 6396 => b"1110101001000",  6397 => b"1110101001000",  6398 => b"1110101000111",  6399 => b"1110101000111",
 6400 => b"1110101000110",  6401 => b"1110101000101",  6402 => b"1110101000101",  6403 => b"1110101000100",
 6404 => b"1110101000011",  6405 => b"1110101000011",  6406 => b"1110101000010",  6407 => b"1110101000001",
 6408 => b"1110101000001",  6409 => b"1110101000000",  6410 => b"1110100111111",  6411 => b"1110100111111",
 6412 => b"1110100111110",  6413 => b"1110100111110",  6414 => b"1110100111101",  6415 => b"1110100111100",
 6416 => b"1110100111100",  6417 => b"1110100111011",  6418 => b"1110100111010",  6419 => b"1110100111010",
 6420 => b"1110100111001",  6421 => b"1110100111000",  6422 => b"1110100111000",  6423 => b"1110100110111",
 6424 => b"1110100110111",  6425 => b"1110100110110",  6426 => b"1110100110101",  6427 => b"1110100110101",
 6428 => b"1110100110100",  6429 => b"1110100110011",  6430 => b"1110100110011",  6431 => b"1110100110010",
 6432 => b"1110100110010",  6433 => b"1110100110001",  6434 => b"1110100110000",  6435 => b"1110100110000",
 6436 => b"1110100101111",  6437 => b"1110100101110",  6438 => b"1110100101110",  6439 => b"1110100101101",
 6440 => b"1110100101101",  6441 => b"1110100101100",  6442 => b"1110100101011",  6443 => b"1110100101011",
 6444 => b"1110100101010",  6445 => b"1110100101010",  6446 => b"1110100101001",  6447 => b"1110100101000",
 6448 => b"1110100101000",  6449 => b"1110100100111",  6450 => b"1110100100110",  6451 => b"1110100100110",
 6452 => b"1110100100101",  6453 => b"1110100100101",  6454 => b"1110100100100",  6455 => b"1110100100011",
 6456 => b"1110100100011",  6457 => b"1110100100010",  6458 => b"1110100100010",  6459 => b"1110100100001",
 6460 => b"1110100100000",  6461 => b"1110100100000",  6462 => b"1110100011111",  6463 => b"1110100011111",
 6464 => b"1110100011110",  6465 => b"1110100011101",  6466 => b"1110100011101",  6467 => b"1110100011100",
 6468 => b"1110100011100",  6469 => b"1110100011011",  6470 => b"1110100011010",  6471 => b"1110100011010",
 6472 => b"1110100011001",  6473 => b"1110100011001",  6474 => b"1110100011000",  6475 => b"1110100011000",
 6476 => b"1110100010111",  6477 => b"1110100010110",  6478 => b"1110100010110",  6479 => b"1110100010101",
 6480 => b"1110100010101",  6481 => b"1110100010100",  6482 => b"1110100010011",  6483 => b"1110100010011",
 6484 => b"1110100010010",  6485 => b"1110100010010",  6486 => b"1110100010001",  6487 => b"1110100010001",
 6488 => b"1110100010000",  6489 => b"1110100001111",  6490 => b"1110100001111",  6491 => b"1110100001110",
 6492 => b"1110100001110",  6493 => b"1110100001101",  6494 => b"1110100001101",  6495 => b"1110100001100",
 6496 => b"1110100001011",  6497 => b"1110100001011",  6498 => b"1110100001010",  6499 => b"1110100001010",
 6500 => b"1110100001001",  6501 => b"1110100001001",  6502 => b"1110100001000",  6503 => b"1110100000111",
 6504 => b"1110100000111",  6505 => b"1110100000110",  6506 => b"1110100000110",  6507 => b"1110100000101",
 6508 => b"1110100000101",  6509 => b"1110100000100",  6510 => b"1110100000100",  6511 => b"1110100000011",
 6512 => b"1110100000010",  6513 => b"1110100000010",  6514 => b"1110100000001",  6515 => b"1110100000001",
 6516 => b"1110100000000",  6517 => b"1110100000000",  6518 => b"1110011111111",  6519 => b"1110011111111",
 6520 => b"1110011111110",  6521 => b"1110011111101",  6522 => b"1110011111101",  6523 => b"1110011111100",
 6524 => b"1110011111100",  6525 => b"1110011111011",  6526 => b"1110011111011",  6527 => b"1110011111010",
 6528 => b"1110011111010",  6529 => b"1110011111001",  6530 => b"1110011111001",  6531 => b"1110011111000",
 6532 => b"1110011111000",  6533 => b"1110011110111",  6534 => b"1110011110110",  6535 => b"1110011110110",
 6536 => b"1110011110101",  6537 => b"1110011110101",  6538 => b"1110011110100",  6539 => b"1110011110100",
 6540 => b"1110011110011",  6541 => b"1110011110011",  6542 => b"1110011110010",  6543 => b"1110011110010",
 6544 => b"1110011110001",  6545 => b"1110011110001",  6546 => b"1110011110000",  6547 => b"1110011110000",
 6548 => b"1110011101111",  6549 => b"1110011101111",  6550 => b"1110011101110",  6551 => b"1110011101110",
 6552 => b"1110011101101",  6553 => b"1110011101101",  6554 => b"1110011101100",  6555 => b"1110011101011",
 6556 => b"1110011101011",  6557 => b"1110011101010",  6558 => b"1110011101010",  6559 => b"1110011101001",
 6560 => b"1110011101001",  6561 => b"1110011101000",  6562 => b"1110011101000",  6563 => b"1110011100111",
 6564 => b"1110011100111",  6565 => b"1110011100110",  6566 => b"1110011100110",  6567 => b"1110011100101",
 6568 => b"1110011100101",  6569 => b"1110011100100",  6570 => b"1110011100100",  6571 => b"1110011100011",
 6572 => b"1110011100011",  6573 => b"1110011100010",  6574 => b"1110011100010",  6575 => b"1110011100001",
 6576 => b"1110011100001",  6577 => b"1110011100000",  6578 => b"1110011100000",  6579 => b"1110011011111",
 6580 => b"1110011011111",  6581 => b"1110011011111",  6582 => b"1110011011110",  6583 => b"1110011011110",
 6584 => b"1110011011101",  6585 => b"1110011011101",  6586 => b"1110011011100",  6587 => b"1110011011100",
 6588 => b"1110011011011",  6589 => b"1110011011011",  6590 => b"1110011011010",  6591 => b"1110011011010",
 6592 => b"1110011011001",  6593 => b"1110011011001",  6594 => b"1110011011000",  6595 => b"1110011011000",
 6596 => b"1110011010111",  6597 => b"1110011010111",  6598 => b"1110011010110",  6599 => b"1110011010110",
 6600 => b"1110011010101",  6601 => b"1110011010101",  6602 => b"1110011010101",  6603 => b"1110011010100",
 6604 => b"1110011010100",  6605 => b"1110011010011",  6606 => b"1110011010011",  6607 => b"1110011010010",
 6608 => b"1110011010010",  6609 => b"1110011010001",  6610 => b"1110011010001",  6611 => b"1110011010000",
 6612 => b"1110011010000",  6613 => b"1110011010000",  6614 => b"1110011001111",  6615 => b"1110011001111",
 6616 => b"1110011001110",  6617 => b"1110011001110",  6618 => b"1110011001101",  6619 => b"1110011001101",
 6620 => b"1110011001100",  6621 => b"1110011001100",  6622 => b"1110011001011",  6623 => b"1110011001011",
 6624 => b"1110011001011",  6625 => b"1110011001010",  6626 => b"1110011001010",  6627 => b"1110011001001",
 6628 => b"1110011001001",  6629 => b"1110011001000",  6630 => b"1110011001000",  6631 => b"1110011001000",
 6632 => b"1110011000111",  6633 => b"1110011000111",  6634 => b"1110011000110",  6635 => b"1110011000110",
 6636 => b"1110011000101",  6637 => b"1110011000101",  6638 => b"1110011000101",  6639 => b"1110011000100",
 6640 => b"1110011000100",  6641 => b"1110011000011",  6642 => b"1110011000011",  6643 => b"1110011000010",
 6644 => b"1110011000010",  6645 => b"1110011000010",  6646 => b"1110011000001",  6647 => b"1110011000001",
 6648 => b"1110011000000",  6649 => b"1110011000000",  6650 => b"1110011000000",  6651 => b"1110010111111",
 6652 => b"1110010111111",  6653 => b"1110010111110",  6654 => b"1110010111110",  6655 => b"1110010111110",
 6656 => b"1110010111101",  6657 => b"1110010111101",  6658 => b"1110010111100",  6659 => b"1110010111100",
 6660 => b"1110010111011",  6661 => b"1110010111011",  6662 => b"1110010111011",  6663 => b"1110010111010",
 6664 => b"1110010111010",  6665 => b"1110010111010",  6666 => b"1110010111001",  6667 => b"1110010111001",
 6668 => b"1110010111000",  6669 => b"1110010111000",  6670 => b"1110010111000",  6671 => b"1110010110111",
 6672 => b"1110010110111",  6673 => b"1110010110110",  6674 => b"1110010110110",  6675 => b"1110010110110",
 6676 => b"1110010110101",  6677 => b"1110010110101",  6678 => b"1110010110100",  6679 => b"1110010110100",
 6680 => b"1110010110100",  6681 => b"1110010110011",  6682 => b"1110010110011",  6683 => b"1110010110011",
 6684 => b"1110010110010",  6685 => b"1110010110010",  6686 => b"1110010110001",  6687 => b"1110010110001",
 6688 => b"1110010110001",  6689 => b"1110010110000",  6690 => b"1110010110000",  6691 => b"1110010110000",
 6692 => b"1110010101111",  6693 => b"1110010101111",  6694 => b"1110010101111",  6695 => b"1110010101110",
 6696 => b"1110010101110",  6697 => b"1110010101101",  6698 => b"1110010101101",  6699 => b"1110010101101",
 6700 => b"1110010101100",  6701 => b"1110010101100",  6702 => b"1110010101100",  6703 => b"1110010101011",
 6704 => b"1110010101011",  6705 => b"1110010101011",  6706 => b"1110010101010",  6707 => b"1110010101010",
 6708 => b"1110010101010",  6709 => b"1110010101001",  6710 => b"1110010101001",  6711 => b"1110010101001",
 6712 => b"1110010101000",  6713 => b"1110010101000",  6714 => b"1110010101000",  6715 => b"1110010100111",
 6716 => b"1110010100111",  6717 => b"1110010100111",  6718 => b"1110010100110",  6719 => b"1110010100110",
 6720 => b"1110010100110",  6721 => b"1110010100101",  6722 => b"1110010100101",  6723 => b"1110010100101",
 6724 => b"1110010100100",  6725 => b"1110010100100",  6726 => b"1110010100100",  6727 => b"1110010100011",
 6728 => b"1110010100011",  6729 => b"1110010100011",  6730 => b"1110010100010",  6731 => b"1110010100010",
 6732 => b"1110010100010",  6733 => b"1110010100001",  6734 => b"1110010100001",  6735 => b"1110010100001",
 6736 => b"1110010100000",  6737 => b"1110010100000",  6738 => b"1110010100000",  6739 => b"1110010100000",
 6740 => b"1110010011111",  6741 => b"1110010011111",  6742 => b"1110010011111",  6743 => b"1110010011110",
 6744 => b"1110010011110",  6745 => b"1110010011110",  6746 => b"1110010011101",  6747 => b"1110010011101",
 6748 => b"1110010011101",  6749 => b"1110010011101",  6750 => b"1110010011100",  6751 => b"1110010011100",
 6752 => b"1110010011100",  6753 => b"1110010011011",  6754 => b"1110010011011",  6755 => b"1110010011011",
 6756 => b"1110010011011",  6757 => b"1110010011010",  6758 => b"1110010011010",  6759 => b"1110010011010",
 6760 => b"1110010011001",  6761 => b"1110010011001",  6762 => b"1110010011001",  6763 => b"1110010011001",
 6764 => b"1110010011000",  6765 => b"1110010011000",  6766 => b"1110010011000",  6767 => b"1110010010111",
 6768 => b"1110010010111",  6769 => b"1110010010111",  6770 => b"1110010010111",  6771 => b"1110010010110",
 6772 => b"1110010010110",  6773 => b"1110010010110",  6774 => b"1110010010110",  6775 => b"1110010010101",
 6776 => b"1110010010101",  6777 => b"1110010010101",  6778 => b"1110010010101",  6779 => b"1110010010100",
 6780 => b"1110010010100",  6781 => b"1110010010100",  6782 => b"1110010010100",  6783 => b"1110010010011",
 6784 => b"1110010010011",  6785 => b"1110010010011",  6786 => b"1110010010011",  6787 => b"1110010010010",
 6788 => b"1110010010010",  6789 => b"1110010010010",  6790 => b"1110010010010",  6791 => b"1110010010001",
 6792 => b"1110010010001",  6793 => b"1110010010001",  6794 => b"1110010010001",  6795 => b"1110010010000",
 6796 => b"1110010010000",  6797 => b"1110010010000",  6798 => b"1110010010000",  6799 => b"1110010001111",
 6800 => b"1110010001111",  6801 => b"1110010001111",  6802 => b"1110010001111",  6803 => b"1110010001111",
 6804 => b"1110010001110",  6805 => b"1110010001110",  6806 => b"1110010001110",  6807 => b"1110010001110",
 6808 => b"1110010001101",  6809 => b"1110010001101",  6810 => b"1110010001101",  6811 => b"1110010001101",
 6812 => b"1110010001101",  6813 => b"1110010001100",  6814 => b"1110010001100",  6815 => b"1110010001100",
 6816 => b"1110010001100",  6817 => b"1110010001011",  6818 => b"1110010001011",  6819 => b"1110010001011",
 6820 => b"1110010001011",  6821 => b"1110010001011",  6822 => b"1110010001010",  6823 => b"1110010001010",
 6824 => b"1110010001010",  6825 => b"1110010001010",  6826 => b"1110010001010",  6827 => b"1110010001001",
 6828 => b"1110010001001",  6829 => b"1110010001001",  6830 => b"1110010001001",  6831 => b"1110010001001",
 6832 => b"1110010001001",  6833 => b"1110010001000",  6834 => b"1110010001000",  6835 => b"1110010001000",
 6836 => b"1110010001000",  6837 => b"1110010001000",  6838 => b"1110010000111",  6839 => b"1110010000111",
 6840 => b"1110010000111",  6841 => b"1110010000111",  6842 => b"1110010000111",  6843 => b"1110010000111",
 6844 => b"1110010000110",  6845 => b"1110010000110",  6846 => b"1110010000110",  6847 => b"1110010000110",
 6848 => b"1110010000110",  6849 => b"1110010000101",  6850 => b"1110010000101",  6851 => b"1110010000101",
 6852 => b"1110010000101",  6853 => b"1110010000101",  6854 => b"1110010000101",  6855 => b"1110010000101",
 6856 => b"1110010000100",  6857 => b"1110010000100",  6858 => b"1110010000100",  6859 => b"1110010000100",
 6860 => b"1110010000100",  6861 => b"1110010000100",  6862 => b"1110010000011",  6863 => b"1110010000011",
 6864 => b"1110010000011",  6865 => b"1110010000011",  6866 => b"1110010000011",  6867 => b"1110010000011",
 6868 => b"1110010000011",  6869 => b"1110010000010",  6870 => b"1110010000010",  6871 => b"1110010000010",
 6872 => b"1110010000010",  6873 => b"1110010000010",  6874 => b"1110010000010",  6875 => b"1110010000010",
 6876 => b"1110010000001",  6877 => b"1110010000001",  6878 => b"1110010000001",  6879 => b"1110010000001",
 6880 => b"1110010000001",  6881 => b"1110010000001",  6882 => b"1110010000001",  6883 => b"1110010000001",
 6884 => b"1110010000000",  6885 => b"1110010000000",  6886 => b"1110010000000",  6887 => b"1110010000000",
 6888 => b"1110010000000",  6889 => b"1110010000000",  6890 => b"1110010000000",  6891 => b"1110010000000",
 6892 => b"1110010000000",  6893 => b"1110001111111",  6894 => b"1110001111111",  6895 => b"1110001111111",
 6896 => b"1110001111111",  6897 => b"1110001111111",  6898 => b"1110001111111",  6899 => b"1110001111111",
 6900 => b"1110001111111",  6901 => b"1110001111111",  6902 => b"1110001111111",  6903 => b"1110001111110",
 6904 => b"1110001111110",  6905 => b"1110001111110",  6906 => b"1110001111110",  6907 => b"1110001111110",
 6908 => b"1110001111110",  6909 => b"1110001111110",  6910 => b"1110001111110",  6911 => b"1110001111110",
 6912 => b"1110001111110",  6913 => b"1110001111110",  6914 => b"1110001111110",  6915 => b"1110001111101",
 6916 => b"1110001111101",  6917 => b"1110001111101",  6918 => b"1110001111101",  6919 => b"1110001111101",
 6920 => b"1110001111101",  6921 => b"1110001111101",  6922 => b"1110001111101",  6923 => b"1110001111101",
 6924 => b"1110001111101",  6925 => b"1110001111101",  6926 => b"1110001111101",  6927 => b"1110001111101",
 6928 => b"1110001111101",  6929 => b"1110001111101",  6930 => b"1110001111100",  6931 => b"1110001111100",
 6932 => b"1110001111100",  6933 => b"1110001111100",  6934 => b"1110001111100",  6935 => b"1110001111100",
 6936 => b"1110001111100",  6937 => b"1110001111100",  6938 => b"1110001111100",  6939 => b"1110001111100",
 6940 => b"1110001111100",  6941 => b"1110001111100",  6942 => b"1110001111100",  6943 => b"1110001111100",
 6944 => b"1110001111100",  6945 => b"1110001111100",  6946 => b"1110001111100",  6947 => b"1110001111100",
 6948 => b"1110001111100",  6949 => b"1110001111100",  6950 => b"1110001111100",  6951 => b"1110001111100",
 6952 => b"1110001111100",  6953 => b"1110001111100",  6954 => b"1110001111011",  6955 => b"1110001111011",
 6956 => b"1110001111011",  6957 => b"1110001111011",  6958 => b"1110001111011",  6959 => b"1110001111011",
 6960 => b"1110001111011",  6961 => b"1110001111011",  6962 => b"1110001111011",  6963 => b"1110001111011",
 6964 => b"1110001111011",  6965 => b"1110001111011",  6966 => b"1110001111011",  6967 => b"1110001111011",
 6968 => b"1110001111011",  6969 => b"1110001111011",  6970 => b"1110001111011",  6971 => b"1110001111011",
 6972 => b"1110001111011",  6973 => b"1110001111011",  6974 => b"1110001111011",  6975 => b"1110001111011",
 6976 => b"1110001111011",  6977 => b"1110001111011",  6978 => b"1110001111011",  6979 => b"1110001111011",
 6980 => b"1110001111011",  6981 => b"1110001111011",  6982 => b"1110001111011",  6983 => b"1110001111011",
 6984 => b"1110001111011",  6985 => b"1110001111011",  6986 => b"1110001111011",  6987 => b"1110001111011",
 6988 => b"1110001111011",  6989 => b"1110001111100",  6990 => b"1110001111100",  6991 => b"1110001111100",
 6992 => b"1110001111100",  6993 => b"1110001111100",  6994 => b"1110001111100",  6995 => b"1110001111100",
 6996 => b"1110001111100",  6997 => b"1110001111100",  6998 => b"1110001111100",  6999 => b"1110001111100",
 7000 => b"1110001111100",  7001 => b"1110001111100",  7002 => b"1110001111100",  7003 => b"1110001111100",
 7004 => b"1110001111100",  7005 => b"1110001111100",  7006 => b"1110001111100",  7007 => b"1110001111100",
 7008 => b"1110001111100",  7009 => b"1110001111100",  7010 => b"1110001111100",  7011 => b"1110001111100",
 7012 => b"1110001111100",  7013 => b"1110001111101",  7014 => b"1110001111101",  7015 => b"1110001111101",
 7016 => b"1110001111101",  7017 => b"1110001111101",  7018 => b"1110001111101",  7019 => b"1110001111101",
 7020 => b"1110001111101",  7021 => b"1110001111101",  7022 => b"1110001111101",  7023 => b"1110001111101",
 7024 => b"1110001111101",  7025 => b"1110001111101",  7026 => b"1110001111101",  7027 => b"1110001111101",
 7028 => b"1110001111110",  7029 => b"1110001111110",  7030 => b"1110001111110",  7031 => b"1110001111110",
 7032 => b"1110001111110",  7033 => b"1110001111110",  7034 => b"1110001111110",  7035 => b"1110001111110",
 7036 => b"1110001111110",  7037 => b"1110001111110",  7038 => b"1110001111110",  7039 => b"1110001111111",
 7040 => b"1110001111111",  7041 => b"1110001111111",  7042 => b"1110001111111",  7043 => b"1110001111111",
 7044 => b"1110001111111",  7045 => b"1110001111111",  7046 => b"1110001111111",  7047 => b"1110001111111",
 7048 => b"1110001111111",  7049 => b"1110010000000",  7050 => b"1110010000000",  7051 => b"1110010000000",
 7052 => b"1110010000000",  7053 => b"1110010000000",  7054 => b"1110010000000",  7055 => b"1110010000000",
 7056 => b"1110010000000",  7057 => b"1110010000000",  7058 => b"1110010000001",  7059 => b"1110010000001",
 7060 => b"1110010000001",  7061 => b"1110010000001",  7062 => b"1110010000001",  7063 => b"1110010000001",
 7064 => b"1110010000001",  7065 => b"1110010000010",  7066 => b"1110010000010",  7067 => b"1110010000010",
 7068 => b"1110010000010",  7069 => b"1110010000010",  7070 => b"1110010000010",  7071 => b"1110010000010",
 7072 => b"1110010000010",  7073 => b"1110010000011",  7074 => b"1110010000011",  7075 => b"1110010000011",
 7076 => b"1110010000011",  7077 => b"1110010000011",  7078 => b"1110010000011",  7079 => b"1110010000100",
 7080 => b"1110010000100",  7081 => b"1110010000100",  7082 => b"1110010000100",  7083 => b"1110010000100",
 7084 => b"1110010000100",  7085 => b"1110010000100",  7086 => b"1110010000101",  7087 => b"1110010000101",
 7088 => b"1110010000101",  7089 => b"1110010000101",  7090 => b"1110010000101",  7091 => b"1110010000101",
 7092 => b"1110010000110",  7093 => b"1110010000110",  7094 => b"1110010000110",  7095 => b"1110010000110",
 7096 => b"1110010000110",  7097 => b"1110010000110",  7098 => b"1110010000111",  7099 => b"1110010000111",
 7100 => b"1110010000111",  7101 => b"1110010000111",  7102 => b"1110010000111",  7103 => b"1110010001000",
 7104 => b"1110010001000",  7105 => b"1110010001000",  7106 => b"1110010001000",  7107 => b"1110010001000",
 7108 => b"1110010001001",  7109 => b"1110010001001",  7110 => b"1110010001001",  7111 => b"1110010001001",
 7112 => b"1110010001001",  7113 => b"1110010001010",  7114 => b"1110010001010",  7115 => b"1110010001010",
 7116 => b"1110010001010",  7117 => b"1110010001010",  7118 => b"1110010001011",  7119 => b"1110010001011",
 7120 => b"1110010001011",  7121 => b"1110010001011",  7122 => b"1110010001011",  7123 => b"1110010001100",
 7124 => b"1110010001100",  7125 => b"1110010001100",  7126 => b"1110010001100",  7127 => b"1110010001100",
 7128 => b"1110010001101",  7129 => b"1110010001101",  7130 => b"1110010001101",  7131 => b"1110010001101",
 7132 => b"1110010001110",  7133 => b"1110010001110",  7134 => b"1110010001110",  7135 => b"1110010001110",
 7136 => b"1110010001111",  7137 => b"1110010001111",  7138 => b"1110010001111",  7139 => b"1110010001111",
 7140 => b"1110010001111",  7141 => b"1110010010000",  7142 => b"1110010010000",  7143 => b"1110010010000",
 7144 => b"1110010010000",  7145 => b"1110010010001",  7146 => b"1110010010001",  7147 => b"1110010010001",
 7148 => b"1110010010001",  7149 => b"1110010010010",  7150 => b"1110010010010",  7151 => b"1110010010010",
 7152 => b"1110010010010",  7153 => b"1110010010011",  7154 => b"1110010010011",  7155 => b"1110010010011",
 7156 => b"1110010010011",  7157 => b"1110010010100",  7158 => b"1110010010100",  7159 => b"1110010010100",
 7160 => b"1110010010101",  7161 => b"1110010010101",  7162 => b"1110010010101",  7163 => b"1110010010101",
 7164 => b"1110010010110",  7165 => b"1110010010110",  7166 => b"1110010010110",  7167 => b"1110010010110",
 7168 => b"1110010010111",  7169 => b"1110010010111",  7170 => b"1110010010111",  7171 => b"1110010011000",
 7172 => b"1110010011000",  7173 => b"1110010011000",  7174 => b"1110010011000",  7175 => b"1110010011001",
 7176 => b"1110010011001",  7177 => b"1110010011001",  7178 => b"1110010011010",  7179 => b"1110010011010",
 7180 => b"1110010011010",  7181 => b"1110010011010",  7182 => b"1110010011011",  7183 => b"1110010011011",
 7184 => b"1110010011011",  7185 => b"1110010011100",  7186 => b"1110010011100",  7187 => b"1110010011100",
 7188 => b"1110010011101",  7189 => b"1110010011101",  7190 => b"1110010011101",  7191 => b"1110010011101",
 7192 => b"1110010011110",  7193 => b"1110010011110",  7194 => b"1110010011110",  7195 => b"1110010011111",
 7196 => b"1110010011111",  7197 => b"1110010011111",  7198 => b"1110010100000",  7199 => b"1110010100000",
 7200 => b"1110010100000",  7201 => b"1110010100001",  7202 => b"1110010100001",  7203 => b"1110010100001",
 7204 => b"1110010100010",  7205 => b"1110010100010",  7206 => b"1110010100010",  7207 => b"1110010100011",
 7208 => b"1110010100011",  7209 => b"1110010100011",  7210 => b"1110010100100",  7211 => b"1110010100100",
 7212 => b"1110010100100",  7213 => b"1110010100101",  7214 => b"1110010100101",  7215 => b"1110010100101",
 7216 => b"1110010100110",  7217 => b"1110010100110",  7218 => b"1110010100110",  7219 => b"1110010100111",
 7220 => b"1110010100111",  7221 => b"1110010100111",  7222 => b"1110010101000",  7223 => b"1110010101000",
 7224 => b"1110010101001",  7225 => b"1110010101001",  7226 => b"1110010101001",  7227 => b"1110010101010",
 7228 => b"1110010101010",  7229 => b"1110010101010",  7230 => b"1110010101011",  7231 => b"1110010101011",
 7232 => b"1110010101011",  7233 => b"1110010101100",  7234 => b"1110010101100",  7235 => b"1110010101101",
 7236 => b"1110010101101",  7237 => b"1110010101101",  7238 => b"1110010101110",  7239 => b"1110010101110",
 7240 => b"1110010101110",  7241 => b"1110010101111",  7242 => b"1110010101111",  7243 => b"1110010110000",
 7244 => b"1110010110000",  7245 => b"1110010110000",  7246 => b"1110010110001",  7247 => b"1110010110001",
 7248 => b"1110010110010",  7249 => b"1110010110010",  7250 => b"1110010110010",  7251 => b"1110010110011",
 7252 => b"1110010110011",  7253 => b"1110010110100",  7254 => b"1110010110100",  7255 => b"1110010110100",
 7256 => b"1110010110101",  7257 => b"1110010110101",  7258 => b"1110010110110",  7259 => b"1110010110110",
 7260 => b"1110010110110",  7261 => b"1110010110111",  7262 => b"1110010110111",  7263 => b"1110010111000",
 7264 => b"1110010111000",  7265 => b"1110010111000",  7266 => b"1110010111001",  7267 => b"1110010111001",
 7268 => b"1110010111010",  7269 => b"1110010111010",  7270 => b"1110010111010",  7271 => b"1110010111011",
 7272 => b"1110010111011",  7273 => b"1110010111100",  7274 => b"1110010111100",  7275 => b"1110010111101",
 7276 => b"1110010111101",  7277 => b"1110010111101",  7278 => b"1110010111110",  7279 => b"1110010111110",
 7280 => b"1110010111111",  7281 => b"1110010111111",  7282 => b"1110011000000",  7283 => b"1110011000000",
 7284 => b"1110011000001",  7285 => b"1110011000001",  7286 => b"1110011000001",  7287 => b"1110011000010",
 7288 => b"1110011000010",  7289 => b"1110011000011",  7290 => b"1110011000011",  7291 => b"1110011000100",
 7292 => b"1110011000100",  7293 => b"1110011000101",  7294 => b"1110011000101",  7295 => b"1110011000101",
 7296 => b"1110011000110",  7297 => b"1110011000110",  7298 => b"1110011000111",  7299 => b"1110011000111",
 7300 => b"1110011001000",  7301 => b"1110011001000",  7302 => b"1110011001001",  7303 => b"1110011001001",
 7304 => b"1110011001010",  7305 => b"1110011001010",  7306 => b"1110011001011",  7307 => b"1110011001011",
 7308 => b"1110011001100",  7309 => b"1110011001100",  7310 => b"1110011001100",  7311 => b"1110011001101",
 7312 => b"1110011001101",  7313 => b"1110011001110",  7314 => b"1110011001110",  7315 => b"1110011001111",
 7316 => b"1110011001111",  7317 => b"1110011010000",  7318 => b"1110011010000",  7319 => b"1110011010001",
 7320 => b"1110011010001",  7321 => b"1110011010010",  7322 => b"1110011010010",  7323 => b"1110011010011",
 7324 => b"1110011010011",  7325 => b"1110011010100",  7326 => b"1110011010100",  7327 => b"1110011010101",
 7328 => b"1110011010101",  7329 => b"1110011010110",  7330 => b"1110011010110",  7331 => b"1110011010111",
 7332 => b"1110011010111",  7333 => b"1110011011000",  7334 => b"1110011011000",  7335 => b"1110011011001",
 7336 => b"1110011011001",  7337 => b"1110011011010",  7338 => b"1110011011010",  7339 => b"1110011011011",
 7340 => b"1110011011011",  7341 => b"1110011011100",  7342 => b"1110011011100",  7343 => b"1110011011101",
 7344 => b"1110011011101",  7345 => b"1110011011110",  7346 => b"1110011011111",  7347 => b"1110011011111",
 7348 => b"1110011100000",  7349 => b"1110011100000",  7350 => b"1110011100001",  7351 => b"1110011100001",
 7352 => b"1110011100010",  7353 => b"1110011100010",  7354 => b"1110011100011",  7355 => b"1110011100011",
 7356 => b"1110011100100",  7357 => b"1110011100100",  7358 => b"1110011100101",  7359 => b"1110011100101",
 7360 => b"1110011100110",  7361 => b"1110011100111",  7362 => b"1110011100111",  7363 => b"1110011101000",
 7364 => b"1110011101000",  7365 => b"1110011101001",  7366 => b"1110011101001",  7367 => b"1110011101010",
 7368 => b"1110011101010",  7369 => b"1110011101011",  7370 => b"1110011101100",  7371 => b"1110011101100",
 7372 => b"1110011101101",  7373 => b"1110011101101",  7374 => b"1110011101110",  7375 => b"1110011101110",
 7376 => b"1110011101111",  7377 => b"1110011101111",  7378 => b"1110011110000",  7379 => b"1110011110001",
 7380 => b"1110011110001",  7381 => b"1110011110010",  7382 => b"1110011110010",  7383 => b"1110011110011",
 7384 => b"1110011110011",  7385 => b"1110011110100",  7386 => b"1110011110101",  7387 => b"1110011110101",
 7388 => b"1110011110110",  7389 => b"1110011110110",  7390 => b"1110011110111",  7391 => b"1110011111000",
 7392 => b"1110011111000",  7393 => b"1110011111001",  7394 => b"1110011111001",  7395 => b"1110011111010",
 7396 => b"1110011111011",  7397 => b"1110011111011",  7398 => b"1110011111100",  7399 => b"1110011111100",
 7400 => b"1110011111101",  7401 => b"1110011111101",  7402 => b"1110011111110",  7403 => b"1110011111111",
 7404 => b"1110011111111",  7405 => b"1110100000000",  7406 => b"1110100000000",  7407 => b"1110100000001",
 7408 => b"1110100000010",  7409 => b"1110100000010",  7410 => b"1110100000011",  7411 => b"1110100000100",
 7412 => b"1110100000100",  7413 => b"1110100000101",  7414 => b"1110100000101",  7415 => b"1110100000110",
 7416 => b"1110100000111",  7417 => b"1110100000111",  7418 => b"1110100001000",  7419 => b"1110100001000",
 7420 => b"1110100001001",  7421 => b"1110100001010",  7422 => b"1110100001010",  7423 => b"1110100001011",
 7424 => b"1110100001100",  7425 => b"1110100001100",  7426 => b"1110100001101",  7427 => b"1110100001101",
 7428 => b"1110100001110",  7429 => b"1110100001111",  7430 => b"1110100001111",  7431 => b"1110100010000",
 7432 => b"1110100010001",  7433 => b"1110100010001",  7434 => b"1110100010010",  7435 => b"1110100010011",
 7436 => b"1110100010011",  7437 => b"1110100010100",  7438 => b"1110100010101",  7439 => b"1110100010101",
 7440 => b"1110100010110",  7441 => b"1110100010110",  7442 => b"1110100010111",  7443 => b"1110100011000",
 7444 => b"1110100011000",  7445 => b"1110100011001",  7446 => b"1110100011010",  7447 => b"1110100011010",
 7448 => b"1110100011011",  7449 => b"1110100011100",  7450 => b"1110100011100",  7451 => b"1110100011101",
 7452 => b"1110100011110",  7453 => b"1110100011110",  7454 => b"1110100011111",  7455 => b"1110100100000",
 7456 => b"1110100100000",  7457 => b"1110100100001",  7458 => b"1110100100010",  7459 => b"1110100100010",
 7460 => b"1110100100011",  7461 => b"1110100100100",  7462 => b"1110100100100",  7463 => b"1110100100101",
 7464 => b"1110100100110",  7465 => b"1110100100110",  7466 => b"1110100100111",  7467 => b"1110100101000",
 7468 => b"1110100101000",  7469 => b"1110100101001",  7470 => b"1110100101010",  7471 => b"1110100101011",
 7472 => b"1110100101011",  7473 => b"1110100101100",  7474 => b"1110100101101",  7475 => b"1110100101101",
 7476 => b"1110100101110",  7477 => b"1110100101111",  7478 => b"1110100101111",  7479 => b"1110100110000",
 7480 => b"1110100110001",  7481 => b"1110100110001",  7482 => b"1110100110010",  7483 => b"1110100110011",
 7484 => b"1110100110100",  7485 => b"1110100110100",  7486 => b"1110100110101",  7487 => b"1110100110110",
 7488 => b"1110100110110",  7489 => b"1110100110111",  7490 => b"1110100111000",  7491 => b"1110100111001",
 7492 => b"1110100111001",  7493 => b"1110100111010",  7494 => b"1110100111011",  7495 => b"1110100111011",
 7496 => b"1110100111100",  7497 => b"1110100111101",  7498 => b"1110100111110",  7499 => b"1110100111110",
 7500 => b"1110100111111",  7501 => b"1110101000000",  7502 => b"1110101000000",  7503 => b"1110101000001",
 7504 => b"1110101000010",  7505 => b"1110101000011",  7506 => b"1110101000011",  7507 => b"1110101000100",
 7508 => b"1110101000101",  7509 => b"1110101000110",  7510 => b"1110101000110",  7511 => b"1110101000111",
 7512 => b"1110101001000",  7513 => b"1110101001000",  7514 => b"1110101001001",  7515 => b"1110101001010",
 7516 => b"1110101001011",  7517 => b"1110101001011",  7518 => b"1110101001100",  7519 => b"1110101001101",
 7520 => b"1110101001110",  7521 => b"1110101001110",  7522 => b"1110101001111",  7523 => b"1110101010000",
 7524 => b"1110101010001",  7525 => b"1110101010001",  7526 => b"1110101010010",  7527 => b"1110101010011",
 7528 => b"1110101010100",  7529 => b"1110101010100",  7530 => b"1110101010101",  7531 => b"1110101010110",
 7532 => b"1110101010111",  7533 => b"1110101010111",  7534 => b"1110101011000",  7535 => b"1110101011001",
 7536 => b"1110101011010",  7537 => b"1110101011011",  7538 => b"1110101011011",  7539 => b"1110101011100",
 7540 => b"1110101011101",  7541 => b"1110101011110",  7542 => b"1110101011110",  7543 => b"1110101011111",
 7544 => b"1110101100000",  7545 => b"1110101100001",  7546 => b"1110101100001",  7547 => b"1110101100010",
 7548 => b"1110101100011",  7549 => b"1110101100100",  7550 => b"1110101100101",  7551 => b"1110101100101",
 7552 => b"1110101100110",  7553 => b"1110101100111",  7554 => b"1110101101000",  7555 => b"1110101101001",
 7556 => b"1110101101001",  7557 => b"1110101101010",  7558 => b"1110101101011",  7559 => b"1110101101100",
 7560 => b"1110101101100",  7561 => b"1110101101101",  7562 => b"1110101101110",  7563 => b"1110101101111",
 7564 => b"1110101110000",  7565 => b"1110101110000",  7566 => b"1110101110001",  7567 => b"1110101110010",
 7568 => b"1110101110011",  7569 => b"1110101110100",  7570 => b"1110101110100",  7571 => b"1110101110101",
 7572 => b"1110101110110",  7573 => b"1110101110111",  7574 => b"1110101111000",  7575 => b"1110101111000",
 7576 => b"1110101111001",  7577 => b"1110101111010",  7578 => b"1110101111011",  7579 => b"1110101111100",
 7580 => b"1110101111101",  7581 => b"1110101111101",  7582 => b"1110101111110",  7583 => b"1110101111111",
 7584 => b"1110110000000",  7585 => b"1110110000001",  7586 => b"1110110000001",  7587 => b"1110110000010",
 7588 => b"1110110000011",  7589 => b"1110110000100",  7590 => b"1110110000101",  7591 => b"1110110000110",
 7592 => b"1110110000110",  7593 => b"1110110000111",  7594 => b"1110110001000",  7595 => b"1110110001001",
 7596 => b"1110110001010",  7597 => b"1110110001011",  7598 => b"1110110001011",  7599 => b"1110110001100",
 7600 => b"1110110001101",  7601 => b"1110110001110",  7602 => b"1110110001111",  7603 => b"1110110010000",
 7604 => b"1110110010000",  7605 => b"1110110010001",  7606 => b"1110110010010",  7607 => b"1110110010011",
 7608 => b"1110110010100",  7609 => b"1110110010101",  7610 => b"1110110010101",  7611 => b"1110110010110",
 7612 => b"1110110010111",  7613 => b"1110110011000",  7614 => b"1110110011001",  7615 => b"1110110011010",
 7616 => b"1110110011011",  7617 => b"1110110011011",  7618 => b"1110110011100",  7619 => b"1110110011101",
 7620 => b"1110110011110",  7621 => b"1110110011111",  7622 => b"1110110100000",  7623 => b"1110110100001",
 7624 => b"1110110100001",  7625 => b"1110110100010",  7626 => b"1110110100011",  7627 => b"1110110100100",
 7628 => b"1110110100101",  7629 => b"1110110100110",  7630 => b"1110110100111",  7631 => b"1110110101000",
 7632 => b"1110110101000",  7633 => b"1110110101001",  7634 => b"1110110101010",  7635 => b"1110110101011",
 7636 => b"1110110101100",  7637 => b"1110110101101",  7638 => b"1110110101110",  7639 => b"1110110101111",
 7640 => b"1110110101111",  7641 => b"1110110110000",  7642 => b"1110110110001",  7643 => b"1110110110010",
 7644 => b"1110110110011",  7645 => b"1110110110100",  7646 => b"1110110110101",  7647 => b"1110110110110",
 7648 => b"1110110110110",  7649 => b"1110110110111",  7650 => b"1110110111000",  7651 => b"1110110111001",
 7652 => b"1110110111010",  7653 => b"1110110111011",  7654 => b"1110110111100",  7655 => b"1110110111101",
 7656 => b"1110110111110",  7657 => b"1110110111111",  7658 => b"1110110111111",  7659 => b"1110111000000",
 7660 => b"1110111000001",  7661 => b"1110111000010",  7662 => b"1110111000011",  7663 => b"1110111000100",
 7664 => b"1110111000101",  7665 => b"1110111000110",  7666 => b"1110111000111",  7667 => b"1110111001000",
 7668 => b"1110111001000",  7669 => b"1110111001001",  7670 => b"1110111001010",  7671 => b"1110111001011",
 7672 => b"1110111001100",  7673 => b"1110111001101",  7674 => b"1110111001110",  7675 => b"1110111001111",
 7676 => b"1110111010000",  7677 => b"1110111010001",  7678 => b"1110111010010",  7679 => b"1110111010010",
 7680 => b"1110111010011",  7681 => b"1110111010100",  7682 => b"1110111010101",  7683 => b"1110111010110",
 7684 => b"1110111010111",  7685 => b"1110111011000",  7686 => b"1110111011001",  7687 => b"1110111011010",
 7688 => b"1110111011011",  7689 => b"1110111011100",  7690 => b"1110111011101",  7691 => b"1110111011110",
 7692 => b"1110111011110",  7693 => b"1110111011111",  7694 => b"1110111100000",  7695 => b"1110111100001",
 7696 => b"1110111100010",  7697 => b"1110111100011",  7698 => b"1110111100100",  7699 => b"1110111100101",
 7700 => b"1110111100110",  7701 => b"1110111100111",  7702 => b"1110111101000",  7703 => b"1110111101001",
 7704 => b"1110111101010",  7705 => b"1110111101011",  7706 => b"1110111101100",  7707 => b"1110111101101",
 7708 => b"1110111101101",  7709 => b"1110111101110",  7710 => b"1110111101111",  7711 => b"1110111110000",
 7712 => b"1110111110001",  7713 => b"1110111110010",  7714 => b"1110111110011",  7715 => b"1110111110100",
 7716 => b"1110111110101",  7717 => b"1110111110110",  7718 => b"1110111110111",  7719 => b"1110111111000",
 7720 => b"1110111111001",  7721 => b"1110111111010",  7722 => b"1110111111011",  7723 => b"1110111111100",
 7724 => b"1110111111101",  7725 => b"1110111111110",  7726 => b"1110111111111",  7727 => b"1111000000000",
 7728 => b"1111000000001",  7729 => b"1111000000010",  7730 => b"1111000000011",  7731 => b"1111000000011",
 7732 => b"1111000000100",  7733 => b"1111000000101",  7734 => b"1111000000110",  7735 => b"1111000000111",
 7736 => b"1111000001000",  7737 => b"1111000001001",  7738 => b"1111000001010",  7739 => b"1111000001011",
 7740 => b"1111000001100",  7741 => b"1111000001101",  7742 => b"1111000001110",  7743 => b"1111000001111",
 7744 => b"1111000010000",  7745 => b"1111000010001",  7746 => b"1111000010010",  7747 => b"1111000010011",
 7748 => b"1111000010100",  7749 => b"1111000010101",  7750 => b"1111000010110",  7751 => b"1111000010111",
 7752 => b"1111000011000",  7753 => b"1111000011001",  7754 => b"1111000011010",  7755 => b"1111000011011",
 7756 => b"1111000011100",  7757 => b"1111000011101",  7758 => b"1111000011110",  7759 => b"1111000011111",
 7760 => b"1111000100000",  7761 => b"1111000100001",  7762 => b"1111000100010",  7763 => b"1111000100011",
 7764 => b"1111000100100",  7765 => b"1111000100101",  7766 => b"1111000100110",  7767 => b"1111000100111",
 7768 => b"1111000101000",  7769 => b"1111000101001",  7770 => b"1111000101010",  7771 => b"1111000101011",
 7772 => b"1111000101100",  7773 => b"1111000101101",  7774 => b"1111000101110",  7775 => b"1111000101111",
 7776 => b"1111000110000",  7777 => b"1111000110001",  7778 => b"1111000110010",  7779 => b"1111000110011",
 7780 => b"1111000110100",  7781 => b"1111000110101",  7782 => b"1111000110110",  7783 => b"1111000110111",
 7784 => b"1111000111000",  7785 => b"1111000111001",  7786 => b"1111000111010",  7787 => b"1111000111011",
 7788 => b"1111000111100",  7789 => b"1111000111101",  7790 => b"1111000111110",  7791 => b"1111000111111",
 7792 => b"1111001000000",  7793 => b"1111001000001",  7794 => b"1111001000010",  7795 => b"1111001000011",
 7796 => b"1111001000100",  7797 => b"1111001000101",  7798 => b"1111001000110",  7799 => b"1111001000111",
 7800 => b"1111001001000",  7801 => b"1111001001001",  7802 => b"1111001001010",  7803 => b"1111001001011",
 7804 => b"1111001001100",  7805 => b"1111001001101",  7806 => b"1111001001110",  7807 => b"1111001001111",
 7808 => b"1111001010000",  7809 => b"1111001010001",  7810 => b"1111001010010",  7811 => b"1111001010011",
 7812 => b"1111001010101",  7813 => b"1111001010110",  7814 => b"1111001010111",  7815 => b"1111001011000",
 7816 => b"1111001011001",  7817 => b"1111001011010",  7818 => b"1111001011011",  7819 => b"1111001011100",
 7820 => b"1111001011101",  7821 => b"1111001011110",  7822 => b"1111001011111",  7823 => b"1111001100000",
 7824 => b"1111001100001",  7825 => b"1111001100010",  7826 => b"1111001100011",  7827 => b"1111001100100",
 7828 => b"1111001100101",  7829 => b"1111001100110",  7830 => b"1111001100111",  7831 => b"1111001101000",
 7832 => b"1111001101001",  7833 => b"1111001101010",  7834 => b"1111001101011",  7835 => b"1111001101100",
 7836 => b"1111001101110",  7837 => b"1111001101111",  7838 => b"1111001110000",  7839 => b"1111001110001",
 7840 => b"1111001110010",  7841 => b"1111001110011",  7842 => b"1111001110100",  7843 => b"1111001110101",
 7844 => b"1111001110110",  7845 => b"1111001110111",  7846 => b"1111001111000",  7847 => b"1111001111001",
 7848 => b"1111001111010",  7849 => b"1111001111011",  7850 => b"1111001111100",  7851 => b"1111001111101",
 7852 => b"1111001111110",  7853 => b"1111001111111",  7854 => b"1111010000001",  7855 => b"1111010000010",
 7856 => b"1111010000011",  7857 => b"1111010000100",  7858 => b"1111010000101",  7859 => b"1111010000110",
 7860 => b"1111010000111",  7861 => b"1111010001000",  7862 => b"1111010001001",  7863 => b"1111010001010",
 7864 => b"1111010001011",  7865 => b"1111010001100",  7866 => b"1111010001101",  7867 => b"1111010001110",
 7868 => b"1111010001111",  7869 => b"1111010010001",  7870 => b"1111010010010",  7871 => b"1111010010011",
 7872 => b"1111010010100",  7873 => b"1111010010101",  7874 => b"1111010010110",  7875 => b"1111010010111",
 7876 => b"1111010011000",  7877 => b"1111010011001",  7878 => b"1111010011010",  7879 => b"1111010011011",
 7880 => b"1111010011100",  7881 => b"1111010011101",  7882 => b"1111010011111",  7883 => b"1111010100000",
 7884 => b"1111010100001",  7885 => b"1111010100010",  7886 => b"1111010100011",  7887 => b"1111010100100",
 7888 => b"1111010100101",  7889 => b"1111010100110",  7890 => b"1111010100111",  7891 => b"1111010101000",
 7892 => b"1111010101001",  7893 => b"1111010101010",  7894 => b"1111010101100",  7895 => b"1111010101101",
 7896 => b"1111010101110",  7897 => b"1111010101111",  7898 => b"1111010110000",  7899 => b"1111010110001",
 7900 => b"1111010110010",  7901 => b"1111010110011",  7902 => b"1111010110100",  7903 => b"1111010110101",
 7904 => b"1111010110110",  7905 => b"1111010111000",  7906 => b"1111010111001",  7907 => b"1111010111010",
 7908 => b"1111010111011",  7909 => b"1111010111100",  7910 => b"1111010111101",  7911 => b"1111010111110",
 7912 => b"1111010111111",  7913 => b"1111011000000",  7914 => b"1111011000001",  7915 => b"1111011000011",
 7916 => b"1111011000100",  7917 => b"1111011000101",  7918 => b"1111011000110",  7919 => b"1111011000111",
 7920 => b"1111011001000",  7921 => b"1111011001001",  7922 => b"1111011001010",  7923 => b"1111011001011",
 7924 => b"1111011001100",  7925 => b"1111011001110",  7926 => b"1111011001111",  7927 => b"1111011010000",
 7928 => b"1111011010001",  7929 => b"1111011010010",  7930 => b"1111011010011",  7931 => b"1111011010100",
 7932 => b"1111011010101",  7933 => b"1111011010110",  7934 => b"1111011011000",  7935 => b"1111011011001",
 7936 => b"1111011011010",  7937 => b"1111011011011",  7938 => b"1111011011100",  7939 => b"1111011011101",
 7940 => b"1111011011110",  7941 => b"1111011011111",  7942 => b"1111011100000",  7943 => b"1111011100010",
 7944 => b"1111011100011",  7945 => b"1111011100100",  7946 => b"1111011100101",  7947 => b"1111011100110",
 7948 => b"1111011100111",  7949 => b"1111011101000",  7950 => b"1111011101001",  7951 => b"1111011101010",
 7952 => b"1111011101100",  7953 => b"1111011101101",  7954 => b"1111011101110",  7955 => b"1111011101111",
 7956 => b"1111011110000",  7957 => b"1111011110001",  7958 => b"1111011110010",  7959 => b"1111011110011",
 7960 => b"1111011110101",  7961 => b"1111011110110",  7962 => b"1111011110111",  7963 => b"1111011111000",
 7964 => b"1111011111001",  7965 => b"1111011111010",  7966 => b"1111011111011",  7967 => b"1111011111100",
 7968 => b"1111011111110",  7969 => b"1111011111111",  7970 => b"1111100000000",  7971 => b"1111100000001",
 7972 => b"1111100000010",  7973 => b"1111100000011",  7974 => b"1111100000100",  7975 => b"1111100000101",
 7976 => b"1111100000111",  7977 => b"1111100001000",  7978 => b"1111100001001",  7979 => b"1111100001010",
 7980 => b"1111100001011",  7981 => b"1111100001100",  7982 => b"1111100001101",  7983 => b"1111100001111",
 7984 => b"1111100010000",  7985 => b"1111100010001",  7986 => b"1111100010010",  7987 => b"1111100010011",
 7988 => b"1111100010100",  7989 => b"1111100010101",  7990 => b"1111100010110",  7991 => b"1111100011000",
 7992 => b"1111100011001",  7993 => b"1111100011010",  7994 => b"1111100011011",  7995 => b"1111100011100",
 7996 => b"1111100011101",  7997 => b"1111100011110",  7998 => b"1111100100000",  7999 => b"1111100100001",
 8000 => b"1111100100010",  8001 => b"1111100100011",  8002 => b"1111100100100",  8003 => b"1111100100101",
 8004 => b"1111100100110",  8005 => b"1111100101000",  8006 => b"1111100101001",  8007 => b"1111100101010",
 8008 => b"1111100101011",  8009 => b"1111100101100",  8010 => b"1111100101101",  8011 => b"1111100101110",
 8012 => b"1111100110000",  8013 => b"1111100110001",  8014 => b"1111100110010",  8015 => b"1111100110011",
 8016 => b"1111100110100",  8017 => b"1111100110101",  8018 => b"1111100110110",  8019 => b"1111100111000",
 8020 => b"1111100111001",  8021 => b"1111100111010",  8022 => b"1111100111011",  8023 => b"1111100111100",
 8024 => b"1111100111101",  8025 => b"1111100111110",  8026 => b"1111101000000",  8027 => b"1111101000001",
 8028 => b"1111101000010",  8029 => b"1111101000011",  8030 => b"1111101000100",  8031 => b"1111101000101",
 8032 => b"1111101000111",  8033 => b"1111101001000",  8034 => b"1111101001001",  8035 => b"1111101001010",
 8036 => b"1111101001011",  8037 => b"1111101001100",  8038 => b"1111101001101",  8039 => b"1111101001111",
 8040 => b"1111101010000",  8041 => b"1111101010001",  8042 => b"1111101010010",  8043 => b"1111101010011",
 8044 => b"1111101010100",  8045 => b"1111101010110",  8046 => b"1111101010111",  8047 => b"1111101011000",
 8048 => b"1111101011001",  8049 => b"1111101011010",  8050 => b"1111101011011",  8051 => b"1111101011100",
 8052 => b"1111101011110",  8053 => b"1111101011111",  8054 => b"1111101100000",  8055 => b"1111101100001",
 8056 => b"1111101100010",  8057 => b"1111101100011",  8058 => b"1111101100101",  8059 => b"1111101100110",
 8060 => b"1111101100111",  8061 => b"1111101101000",  8062 => b"1111101101001",  8063 => b"1111101101010",
 8064 => b"1111101101100",  8065 => b"1111101101101",  8066 => b"1111101101110",  8067 => b"1111101101111",
 8068 => b"1111101110000",  8069 => b"1111101110001",  8070 => b"1111101110011",  8071 => b"1111101110100",
 8072 => b"1111101110101",  8073 => b"1111101110110",  8074 => b"1111101110111",  8075 => b"1111101111000",
 8076 => b"1111101111010",  8077 => b"1111101111011",  8078 => b"1111101111100",  8079 => b"1111101111101",
 8080 => b"1111101111110",  8081 => b"1111101111111",  8082 => b"1111110000001",  8083 => b"1111110000010",
 8084 => b"1111110000011",  8085 => b"1111110000100",  8086 => b"1111110000101",  8087 => b"1111110000110",
 8088 => b"1111110001000",  8089 => b"1111110001001",  8090 => b"1111110001010",  8091 => b"1111110001011",
 8092 => b"1111110001100",  8093 => b"1111110001101",  8094 => b"1111110001111",  8095 => b"1111110010000",
 8096 => b"1111110010001",  8097 => b"1111110010010",  8098 => b"1111110010011",  8099 => b"1111110010100",
 8100 => b"1111110010110",  8101 => b"1111110010111",  8102 => b"1111110011000",  8103 => b"1111110011001",
 8104 => b"1111110011010",  8105 => b"1111110011011",  8106 => b"1111110011101",  8107 => b"1111110011110",
 8108 => b"1111110011111",  8109 => b"1111110100000",  8110 => b"1111110100001",  8111 => b"1111110100010",
 8112 => b"1111110100100",  8113 => b"1111110100101",  8114 => b"1111110100110",  8115 => b"1111110100111",
 8116 => b"1111110101000",  8117 => b"1111110101001",  8118 => b"1111110101011",  8119 => b"1111110101100",
 8120 => b"1111110101101",  8121 => b"1111110101110",  8122 => b"1111110101111",  8123 => b"1111110110000",
 8124 => b"1111110110010",  8125 => b"1111110110011",  8126 => b"1111110110100",  8127 => b"1111110110101",
 8128 => b"1111110110110",  8129 => b"1111110111000",  8130 => b"1111110111001",  8131 => b"1111110111010",
 8132 => b"1111110111011",  8133 => b"1111110111100",  8134 => b"1111110111101",  8135 => b"1111110111111",
 8136 => b"1111111000000",  8137 => b"1111111000001",  8138 => b"1111111000010",  8139 => b"1111111000011",
 8140 => b"1111111000100",  8141 => b"1111111000110",  8142 => b"1111111000111",  8143 => b"1111111001000",
 8144 => b"1111111001001",  8145 => b"1111111001010",  8146 => b"1111111001100",  8147 => b"1111111001101",
 8148 => b"1111111001110",  8149 => b"1111111001111",  8150 => b"1111111010000",  8151 => b"1111111010001",
 8152 => b"1111111010011",  8153 => b"1111111010100",  8154 => b"1111111010101",  8155 => b"1111111010110",
 8156 => b"1111111010111",  8157 => b"1111111011000",  8158 => b"1111111011010",  8159 => b"1111111011011",
 8160 => b"1111111011100",  8161 => b"1111111011101",  8162 => b"1111111011110",  8163 => b"1111111100000",
 8164 => b"1111111100001",  8165 => b"1111111100010",  8166 => b"1111111100011",  8167 => b"1111111100100",
 8168 => b"1111111100101",  8169 => b"1111111100111",  8170 => b"1111111101000",  8171 => b"1111111101001",
 8172 => b"1111111101010",  8173 => b"1111111101011",  8174 => b"1111111101100",  8175 => b"1111111101110",
 8176 => b"1111111101111",  8177 => b"1111111110000",  8178 => b"1111111110001",  8179 => b"1111111110010",
 8180 => b"1111111110100",  8181 => b"1111111110101",  8182 => b"1111111110110",  8183 => b"1111111110111",
 8184 => b"1111111111000",  8185 => b"1111111111001",  8186 => b"1111111111011",  8187 => b"1111111111100",
 8188 => b"1111111111101",  8189 => b"1111111111110",  8190 => b"1111111111111",  8191 => b"0000000000000" 

);

signal state, nx_state : estado;

signal data_valid : std_logic;

begin

    update_state : process(clk, nrst)
    begin
        if rising_edge(clk) then
            if nrst = '0' then
                state <= init;
            else
                state <= nx_state;
            end if;
        end if;
    end process update_state;


    next_state : process(state)
    begin
        case state is
        when init =>
            n <= 0;
            axis_mtr_tdata <= my_data(n);
            axis_mtr_tvalid <= '0';
            nx_state <= tvalid;
        when tvalid =>
            axis_mtr_tdata <= my_data(n);
            axis_mtr_tvalid <= '1';
            if axis_mtr_tready = '1' then
                nx_state <= tready;
            end if;
        when tready =>
            n <= n+1;
            if n=8191 then n <= 0; end if; -- counter reset at 8191
            axis_mtr_tvalid <= '0';
            nx_state <= tvalid;
        when others =>
            n <= 0;
            axis_mtr_tvalid <= '0';
            axis_mtr_tdata <= my_data(n);
            nx_state <= init;
        end case;
    end process next_state;

end Behavioral;

